// Benchmark "top" written by ABC on Tue Jul 22 21:34:14 2025

module top ( 
    \priority0 , \priority1 , \priority2 , \priority3 ,
    \priority4 , \priority5 , \priority6 , \priority7 ,
    \priority8 , \priority9 , \priority10 , \priority11 ,
    \priority12 , \priority13 , \priority14 , \priority15 ,
    \priority16 , \priority17 , \priority18 , \priority19 ,
    \priority20 , \priority21 , \priority22 , \priority23 ,
    \priority24 , \priority25 , \priority26 , \priority27 ,
    \priority28 , \priority29 , \priority30 , \priority31 ,
    \priority32 , \priority33 , \priority34 , \priority35 ,
    \priority36 , \priority37 , \priority38 , \priority39 ,
    \priority40 , \priority41 , \priority42 , \priority43 ,
    \priority44 , \priority45 , \priority46 , \priority47 ,
    \priority48 , \priority49 , \priority50 , \priority51 ,
    \priority52 , \priority53 , \priority54 , \priority55 ,
    \priority56 , \priority57 , \priority58 , \priority59 ,
    \priority60 , \priority61 , \priority62 , \priority63 ,
    \priority64 , \priority65 , \priority66 , \priority67 ,
    \priority68 , \priority69 , \priority70 , \priority71 ,
    \priority72 , \priority73 , \priority74 , \priority75 ,
    \priority76 , \priority77 , \priority78 , \priority79 ,
    \priority80 , \priority81 , \priority82 , \priority83 ,
    \priority84 , \priority85 , \priority86 , \priority87 ,
    \priority88 , \priority89 , \priority90 , \priority91 ,
    \priority92 , \priority93 , \priority94 , \priority95 ,
    \priority96 , \priority97 , \priority98 , \priority99 ,
    \priority100 , \priority101 , \priority102 , \priority103 ,
    \priority104 , \priority105 , \priority106 , \priority107 ,
    \priority108 , \priority109 , \priority110 , \priority111 ,
    \priority112 , \priority113 , \priority114 , \priority115 ,
    \priority116 , \priority117 , \priority118 , \priority119 ,
    \priority120 , \priority121 , \priority122 , \priority123 ,
    \priority124 , \priority125 , \priority126 , \priority127 ,
    \req0 , \req1 , \req2 , \req3 , \req4 , \req5 , \req6 ,
    \req7 , \req8 , \req9 , \req10 , \req11 , \req12 ,
    \req13 , \req14 , \req15 , \req16 , \req17 , \req18 ,
    \req19 , \req20 , \req21 , \req22 , \req23 , \req24 ,
    \req25 , \req26 , \req27 , \req28 , \req29 , \req30 ,
    \req31 , \req32 , \req33 , \req34 , \req35 , \req36 ,
    \req37 , \req38 , \req39 , \req40 , \req41 , \req42 ,
    \req43 , \req44 , \req45 , \req46 , \req47 , \req48 ,
    \req49 , \req50 , \req51 , \req52 , \req53 , \req54 ,
    \req55 , \req56 , \req57 , \req58 , \req59 , \req60 ,
    \req61 , \req62 , \req63 , \req64 , \req65 , \req66 ,
    \req67 , \req68 , \req69 , \req70 , \req71 , \req72 ,
    \req73 , \req74 , \req75 , \req76 , \req77 , \req78 ,
    \req79 , \req80 , \req81 , \req82 , \req83 , \req84 ,
    \req85 , \req86 , \req87 , \req88 , \req89 , \req90 ,
    \req91 , \req92 , \req93 , \req94 , \req95 , \req96 ,
    \req97 , \req98 , \req99 , \req100 , \req101 , \req102 ,
    \req103 , \req104 , \req105 , \req106 , \req107 , \req108 ,
    \req109 , \req110 , \req111 , \req112 , \req113 , \req114 ,
    \req115 , \req116 , \req117 , \req118 , \req119 , \req120 ,
    \req121 , \req122 , \req123 , \req124 , \req125 , \req126 ,
    \req127 ,
    \grant0 , \grant1 , \grant2 , \grant3 , \grant4 , \grant5 ,
    \grant6 , \grant7 , \grant8 , \grant9 , \grant10 ,
    \grant11 , \grant12 , \grant13 , \grant14 , \grant15 ,
    \grant16 , \grant17 , \grant18 , \grant19 , \grant20 ,
    \grant21 , \grant22 , \grant23 , \grant24 , \grant25 ,
    \grant26 , \grant27 , \grant28 , \grant29 , \grant30 ,
    \grant31 , \grant32 , \grant33 , \grant34 , \grant35 ,
    \grant36 , \grant37 , \grant38 , \grant39 , \grant40 ,
    \grant41 , \grant42 , \grant43 , \grant44 , \grant45 ,
    \grant46 , \grant47 , \grant48 , \grant49 , \grant50 ,
    \grant51 , \grant52 , \grant53 , \grant54 , \grant55 ,
    \grant56 , \grant57 , \grant58 , \grant59 , \grant60 ,
    \grant61 , \grant62 , \grant63 , \grant64 , \grant65 ,
    \grant66 , \grant67 , \grant68 , \grant69 , \grant70 ,
    \grant71 , \grant72 , \grant73 , \grant74 , \grant75 ,
    \grant76 , \grant77 , \grant78 , \grant79 , \grant80 ,
    \grant81 , \grant82 , \grant83 , \grant84 , \grant85 ,
    \grant86 , \grant87 , \grant88 , \grant89 , \grant90 ,
    \grant91 , \grant92 , \grant93 , \grant94 , \grant95 ,
    \grant96 , \grant97 , \grant98 , \grant99 , \grant100 ,
    \grant101 , \grant102 , \grant103 , \grant104 , \grant105 ,
    \grant106 , \grant107 , \grant108 , \grant109 , \grant110 ,
    \grant111 , \grant112 , \grant113 , \grant114 , \grant115 ,
    \grant116 , \grant117 , \grant118 , \grant119 , \grant120 ,
    \grant121 , \grant122 , \grant123 , \grant124 , \grant125 ,
    \grant126 , \grant127 , anyGrant  );
  input  \priority0 , \priority1 , \priority2 , \priority3 ,
    \priority4 , \priority5 , \priority6 , \priority7 ,
    \priority8 , \priority9 , \priority10 , \priority11 ,
    \priority12 , \priority13 , \priority14 , \priority15 ,
    \priority16 , \priority17 , \priority18 , \priority19 ,
    \priority20 , \priority21 , \priority22 , \priority23 ,
    \priority24 , \priority25 , \priority26 , \priority27 ,
    \priority28 , \priority29 , \priority30 , \priority31 ,
    \priority32 , \priority33 , \priority34 , \priority35 ,
    \priority36 , \priority37 , \priority38 , \priority39 ,
    \priority40 , \priority41 , \priority42 , \priority43 ,
    \priority44 , \priority45 , \priority46 , \priority47 ,
    \priority48 , \priority49 , \priority50 , \priority51 ,
    \priority52 , \priority53 , \priority54 , \priority55 ,
    \priority56 , \priority57 , \priority58 , \priority59 ,
    \priority60 , \priority61 , \priority62 , \priority63 ,
    \priority64 , \priority65 , \priority66 , \priority67 ,
    \priority68 , \priority69 , \priority70 , \priority71 ,
    \priority72 , \priority73 , \priority74 , \priority75 ,
    \priority76 , \priority77 , \priority78 , \priority79 ,
    \priority80 , \priority81 , \priority82 , \priority83 ,
    \priority84 , \priority85 , \priority86 , \priority87 ,
    \priority88 , \priority89 , \priority90 , \priority91 ,
    \priority92 , \priority93 , \priority94 , \priority95 ,
    \priority96 , \priority97 , \priority98 , \priority99 ,
    \priority100 , \priority101 , \priority102 , \priority103 ,
    \priority104 , \priority105 , \priority106 , \priority107 ,
    \priority108 , \priority109 , \priority110 , \priority111 ,
    \priority112 , \priority113 , \priority114 , \priority115 ,
    \priority116 , \priority117 , \priority118 , \priority119 ,
    \priority120 , \priority121 , \priority122 , \priority123 ,
    \priority124 , \priority125 , \priority126 , \priority127 ,
    \req0 , \req1 , \req2 , \req3 , \req4 , \req5 , \req6 ,
    \req7 , \req8 , \req9 , \req10 , \req11 , \req12 ,
    \req13 , \req14 , \req15 , \req16 , \req17 , \req18 ,
    \req19 , \req20 , \req21 , \req22 , \req23 , \req24 ,
    \req25 , \req26 , \req27 , \req28 , \req29 , \req30 ,
    \req31 , \req32 , \req33 , \req34 , \req35 , \req36 ,
    \req37 , \req38 , \req39 , \req40 , \req41 , \req42 ,
    \req43 , \req44 , \req45 , \req46 , \req47 , \req48 ,
    \req49 , \req50 , \req51 , \req52 , \req53 , \req54 ,
    \req55 , \req56 , \req57 , \req58 , \req59 , \req60 ,
    \req61 , \req62 , \req63 , \req64 , \req65 , \req66 ,
    \req67 , \req68 , \req69 , \req70 , \req71 , \req72 ,
    \req73 , \req74 , \req75 , \req76 , \req77 , \req78 ,
    \req79 , \req80 , \req81 , \req82 , \req83 , \req84 ,
    \req85 , \req86 , \req87 , \req88 , \req89 , \req90 ,
    \req91 , \req92 , \req93 , \req94 , \req95 , \req96 ,
    \req97 , \req98 , \req99 , \req100 , \req101 , \req102 ,
    \req103 , \req104 , \req105 , \req106 , \req107 , \req108 ,
    \req109 , \req110 , \req111 , \req112 , \req113 , \req114 ,
    \req115 , \req116 , \req117 , \req118 , \req119 , \req120 ,
    \req121 , \req122 , \req123 , \req124 , \req125 , \req126 ,
    \req127 ;
  output \grant0 , \grant1 , \grant2 , \grant3 , \grant4 ,
    \grant5 , \grant6 , \grant7 , \grant8 , \grant9 ,
    \grant10 , \grant11 , \grant12 , \grant13 , \grant14 ,
    \grant15 , \grant16 , \grant17 , \grant18 , \grant19 ,
    \grant20 , \grant21 , \grant22 , \grant23 , \grant24 ,
    \grant25 , \grant26 , \grant27 , \grant28 , \grant29 ,
    \grant30 , \grant31 , \grant32 , \grant33 , \grant34 ,
    \grant35 , \grant36 , \grant37 , \grant38 , \grant39 ,
    \grant40 , \grant41 , \grant42 , \grant43 , \grant44 ,
    \grant45 , \grant46 , \grant47 , \grant48 , \grant49 ,
    \grant50 , \grant51 , \grant52 , \grant53 , \grant54 ,
    \grant55 , \grant56 , \grant57 , \grant58 , \grant59 ,
    \grant60 , \grant61 , \grant62 , \grant63 , \grant64 ,
    \grant65 , \grant66 , \grant67 , \grant68 , \grant69 ,
    \grant70 , \grant71 , \grant72 , \grant73 , \grant74 ,
    \grant75 , \grant76 , \grant77 , \grant78 , \grant79 ,
    \grant80 , \grant81 , \grant82 , \grant83 , \grant84 ,
    \grant85 , \grant86 , \grant87 , \grant88 , \grant89 ,
    \grant90 , \grant91 , \grant92 , \grant93 , \grant94 ,
    \grant95 , \grant96 , \grant97 , \grant98 , \grant99 ,
    \grant100 , \grant101 , \grant102 , \grant103 , \grant104 ,
    \grant105 , \grant106 , \grant107 , \grant108 , \grant109 ,
    \grant110 , \grant111 , \grant112 , \grant113 , \grant114 ,
    \grant115 , \grant116 , \grant117 , \grant118 , \grant119 ,
    \grant120 , \grant121 , \grant122 , \grant123 , \grant124 ,
    \grant125 , \grant126 , \grant127 , anyGrant;
  wire new_n386, new_n387, new_n388, new_n389, new_n390, new_n391, new_n392,
    new_n393, new_n394, new_n395, new_n396, new_n397, new_n398, new_n399,
    new_n400, new_n401, new_n402, new_n403, new_n404, new_n405, new_n406,
    new_n407, new_n408, new_n409, new_n410, new_n411, new_n412, new_n413,
    new_n414, new_n415, new_n416, new_n417, new_n418, new_n419, new_n420,
    new_n421, new_n422, new_n423, new_n424, new_n425, new_n426, new_n427,
    new_n428, new_n429, new_n430, new_n431, new_n432, new_n433, new_n434,
    new_n435, new_n436, new_n437, new_n438, new_n439, new_n440, new_n441,
    new_n442, new_n443, new_n444, new_n445, new_n446, new_n447, new_n448,
    new_n449, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n461, new_n462,
    new_n463, new_n464, new_n465, new_n466, new_n467, new_n468, new_n469,
    new_n470, new_n471, new_n472, new_n473, new_n474, new_n475, new_n476,
    new_n477, new_n478, new_n479, new_n480, new_n481, new_n482, new_n483,
    new_n484, new_n485, new_n486, new_n487, new_n488, new_n489, new_n490,
    new_n491, new_n492, new_n493, new_n494, new_n495, new_n496, new_n497,
    new_n498, new_n499, new_n500, new_n501, new_n502, new_n503, new_n504,
    new_n505, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1033, new_n1034,
    new_n1036, new_n1037, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1051, new_n1052, new_n1053, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1081, new_n1082, new_n1083, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1092,
    new_n1093, new_n1094, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1102, new_n1103, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1115,
    new_n1116, new_n1118, new_n1119, new_n1120, new_n1122, new_n1123,
    new_n1124, new_n1126, new_n1127, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1141, new_n1142, new_n1144, new_n1145, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1160, new_n1161, new_n1162, new_n1164,
    new_n1165, new_n1167, new_n1168, new_n1169, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1190, new_n1191, new_n1192, new_n1193, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1200, new_n1201, new_n1202,
    new_n1204, new_n1205, new_n1206, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1220, new_n1221, new_n1222, new_n1224, new_n1225, new_n1226,
    new_n1228, new_n1229, new_n1230, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1245, new_n1246, new_n1248, new_n1250, new_n1251,
    new_n1252, new_n1254, new_n1255, new_n1256, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1265, new_n1266, new_n1268,
    new_n1269, new_n1270, new_n1272, new_n1273, new_n1274, new_n1276,
    new_n1277, new_n1278, new_n1280, new_n1281, new_n1283, new_n1285,
    new_n1286, new_n1287, new_n1289, new_n1290, new_n1291, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1298, new_n1299, new_n1301,
    new_n1302, new_n1304, new_n1305, new_n1306, new_n1308, new_n1309,
    new_n1310, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1320, new_n1321, new_n1322, new_n1324, new_n1325,
    new_n1326, new_n1328, new_n1329, new_n1331, new_n1332, new_n1333,
    new_n1334, new_n1335, new_n1336, new_n1337, new_n1338, new_n1339,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346, new_n1347,
    new_n1349, new_n1350, new_n1351, new_n1353, new_n1354, new_n1355,
    new_n1356, new_n1358, new_n1359, new_n1360, new_n1361, new_n1363,
    new_n1364, new_n1365, new_n1366, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1377,
    new_n1378, new_n1380, new_n1381, new_n1383, new_n1384, new_n1386,
    new_n1387, new_n1389, new_n1390, new_n1392, new_n1395, new_n1398,
    new_n1399, new_n1401, new_n1402, new_n1403, new_n1405, new_n1407,
    new_n1408, new_n1410, new_n1411, new_n1414, new_n1415, new_n1416,
    new_n1418, new_n1420, new_n1422, new_n1423, new_n1424, new_n1425,
    new_n1426, new_n1427, new_n1428, new_n1429, new_n1430, new_n1431,
    new_n1432, new_n1433, new_n1434, new_n1435, new_n1436, new_n1437,
    new_n1438, new_n1439, new_n1440, new_n1441, new_n1442, new_n1443,
    new_n1444, new_n1445, new_n1446, new_n1447, new_n1448, new_n1449,
    new_n1450, new_n1451, new_n1452, new_n1453, new_n1454, new_n1455,
    new_n1456, new_n1457, new_n1458, new_n1459, new_n1460, new_n1461,
    new_n1462, new_n1463, new_n1464;
  inv1  g0000(.a(\req0 ), .O(new_n386));
  inv1  g0001(.a(\priority121 ), .O(new_n387));
  inv1  g0002(.a(\priority114 ), .O(new_n388));
  inv1  g0003(.a(\priority112 ), .O(new_n389));
  inv1  g0004(.a(\req99 ), .O(new_n390));
  inv1  g0005(.a(\priority97 ), .O(new_n391));
  inv1  g0006(.a(\req93 ), .O(new_n392));
  aoi21 g0007(.a(new_n392), .b(\priority93 ), .c(\priority94 ), .O(new_n393));
  inv1  g0008(.a(\req89 ), .O(new_n394));
  inv1  g0009(.a(\req88 ), .O(new_n395));
  aoi21 g0010(.a(new_n395), .b(\priority88 ), .c(\priority89 ), .O(new_n396));
  inv1  g0011(.a(new_n396), .O(new_n397));
  inv1  g0012(.a(\priority87 ), .O(new_n398));
  inv1  g0013(.a(\req83 ), .O(new_n399));
  aoi21 g0014(.a(new_n399), .b(\priority83 ), .c(\priority84 ), .O(new_n400));
  inv1  g0015(.a(\req79 ), .O(new_n401));
  inv1  g0016(.a(\req78 ), .O(new_n402));
  aoi21 g0017(.a(new_n402), .b(\priority78 ), .c(\priority79 ), .O(new_n403));
  inv1  g0018(.a(new_n403), .O(new_n404));
  inv1  g0019(.a(\priority77 ), .O(new_n405));
  inv1  g0020(.a(\req63 ), .O(new_n406));
  inv1  g0021(.a(\req64 ), .O(new_n407));
  nor2  g0022(.a(\req62 ), .b(\req61 ), .O(new_n408));
  nor2  g0023(.a(\req66 ), .b(\req65 ), .O(new_n409));
  nand4 g0024(.a(new_n409), .b(new_n408), .c(new_n407), .d(new_n406), .O(new_n410));
  inv1  g0025(.a(\req67 ), .O(new_n411));
  inv1  g0026(.a(\req68 ), .O(new_n412));
  nor3  g0027(.a(\req73 ), .b(\req72 ), .c(\req71 ), .O(new_n413));
  nor2  g0028(.a(\req70 ), .b(\req69 ), .O(new_n414));
  nand4 g0029(.a(new_n414), .b(new_n413), .c(new_n412), .d(new_n411), .O(new_n415));
  nor2  g0030(.a(new_n415), .b(new_n410), .O(new_n416));
  inv1  g0031(.a(new_n416), .O(new_n417));
  inv1  g0032(.a(\priority56 ), .O(new_n418));
  inv1  g0033(.a(\req53 ), .O(new_n419));
  inv1  g0034(.a(\priority46 ), .O(new_n420));
  inv1  g0035(.a(\req43 ), .O(new_n421));
  inv1  g0036(.a(\priority36 ), .O(new_n422));
  inv1  g0037(.a(\priority29 ), .O(new_n423));
  inv1  g0038(.a(\req26 ), .O(new_n424));
  inv1  g0039(.a(\priority19 ), .O(new_n425));
  inv1  g0040(.a(\req11 ), .O(new_n426));
  inv1  g0041(.a(\priority4 ), .O(new_n427));
  inv1  g0042(.a(\req1 ), .O(new_n428));
  inv1  g0043(.a(\req121 ), .O(new_n429));
  inv1  g0044(.a(\req122 ), .O(new_n430));
  nor2  g0045(.a(\req120 ), .b(\req119 ), .O(new_n431));
  nor2  g0046(.a(\req124 ), .b(\req123 ), .O(new_n432));
  nand4 g0047(.a(new_n432), .b(new_n431), .c(new_n430), .d(new_n429), .O(new_n433));
  inv1  g0048(.a(new_n433), .O(new_n434));
  inv1  g0049(.a(\req117 ), .O(new_n435));
  inv1  g0050(.a(\priority116 ), .O(new_n436));
  inv1  g0051(.a(\req116 ), .O(new_n437));
  nor2  g0052(.a(\req115 ), .b(\priority117 ), .O(new_n438));
  nand4 g0053(.a(new_n438), .b(new_n437), .c(new_n436), .d(\priority115 ), .O(new_n439));
  aoi21 g0054(.a(new_n437), .b(\priority116 ), .c(\priority117 ), .O(new_n440));
  nand2 g0055(.a(new_n440), .b(new_n439), .O(new_n441));
  nand2 g0056(.a(new_n441), .b(new_n435), .O(new_n442));
  nor2  g0057(.a(\req115 ), .b(\req114 ), .O(new_n443));
  nor2  g0058(.a(\req126 ), .b(\req118 ), .O(new_n444));
  nand4 g0059(.a(new_n444), .b(new_n443), .c(new_n435), .d(new_n437), .O(new_n445));
  inv1  g0060(.a(new_n445), .O(new_n446));
  inv1  g0061(.a(\req113 ), .O(new_n447));
  aoi21 g0062(.a(new_n447), .b(\priority113 ), .c(\priority114 ), .O(new_n448));
  inv1  g0063(.a(\priority113 ), .O(new_n449));
  inv1  g0064(.a(\req112 ), .O(new_n450));
  nor2  g0065(.a(\req113 ), .b(\priority114 ), .O(new_n451));
  nand4 g0066(.a(new_n451), .b(new_n450), .c(new_n449), .d(\priority112 ), .O(new_n452));
  nand2 g0067(.a(new_n452), .b(new_n448), .O(new_n453));
  nand2 g0068(.a(new_n453), .b(new_n446), .O(new_n454));
  inv1  g0069(.a(\priority118 ), .O(new_n455));
  inv1  g0070(.a(\priority119 ), .O(new_n456));
  inv1  g0071(.a(\req118 ), .O(new_n457));
  nand3 g0072(.a(new_n457), .b(new_n456), .c(new_n455), .O(new_n458));
  nor2  g0073(.a(new_n458), .b(new_n433), .O(new_n459));
  nand3 g0074(.a(new_n459), .b(new_n454), .c(new_n442), .O(new_n460));
  nor2  g0075(.a(new_n457), .b(\priority119 ), .O(new_n461));
  nand3 g0076(.a(new_n461), .b(new_n434), .c(new_n454), .O(new_n462));
  nand3 g0077(.a(new_n462), .b(new_n460), .c(new_n434), .O(new_n463));
  nor2  g0078(.a(\req120 ), .b(\priority122 ), .O(new_n464));
  nand4 g0079(.a(new_n464), .b(new_n429), .c(new_n387), .d(\priority120 ), .O(new_n465));
  aoi21 g0080(.a(new_n429), .b(\priority121 ), .c(\priority122 ), .O(new_n466));
  aoi21 g0081(.a(new_n466), .b(new_n465), .c(\req122 ), .O(new_n467));
  inv1  g0082(.a(\priority123 ), .O(new_n468));
  inv1  g0083(.a(\priority124 ), .O(new_n469));
  nand3 g0084(.a(new_n432), .b(new_n469), .c(new_n468), .O(new_n470));
  aoi21 g0085(.a(\req123 ), .b(new_n469), .c(\req124 ), .O(new_n471));
  oai21 g0086(.a(new_n470), .b(new_n467), .c(new_n471), .O(new_n472));
  inv1  g0087(.a(\priority125 ), .O(new_n473));
  inv1  g0088(.a(\priority126 ), .O(new_n474));
  inv1  g0089(.a(\req125 ), .O(new_n475));
  inv1  g0090(.a(\req126 ), .O(new_n476));
  nand4 g0091(.a(new_n476), .b(new_n475), .c(new_n474), .d(new_n473), .O(new_n477));
  inv1  g0092(.a(new_n477), .O(new_n478));
  nand3 g0093(.a(new_n478), .b(new_n472), .c(new_n463), .O(new_n479));
  aoi21 g0094(.a(\req125 ), .b(new_n474), .c(\req126 ), .O(new_n480));
  aoi21 g0095(.a(new_n480), .b(new_n479), .c(\priority127 ), .O(new_n481));
  nor2  g0096(.a(\priority1 ), .b(\priority0 ), .O(new_n482));
  nor2  g0097(.a(\req127 ), .b(\req0 ), .O(new_n483));
  nand2 g0098(.a(new_n483), .b(new_n482), .O(new_n484));
  aoi21 g0099(.a(new_n386), .b(\priority0 ), .c(\priority1 ), .O(new_n485));
  oai21 g0100(.a(new_n484), .b(new_n481), .c(new_n485), .O(new_n486));
  inv1  g0101(.a(\priority2 ), .O(new_n487));
  inv1  g0102(.a(\priority3 ), .O(new_n488));
  inv1  g0103(.a(\req2 ), .O(new_n489));
  inv1  g0104(.a(\req3 ), .O(new_n490));
  nand4 g0105(.a(new_n490), .b(new_n489), .c(new_n488), .d(new_n487), .O(new_n491));
  aoi21 g0106(.a(new_n486), .b(new_n428), .c(new_n491), .O(new_n492));
  oai21 g0107(.a(new_n489), .b(\priority3 ), .c(new_n490), .O(new_n493));
  oai21 g0108(.a(new_n493), .b(new_n492), .c(new_n427), .O(new_n494));
  inv1  g0109(.a(\priority5 ), .O(new_n495));
  inv1  g0110(.a(\priority6 ), .O(new_n496));
  inv1  g0111(.a(\req4 ), .O(new_n497));
  inv1  g0112(.a(\req5 ), .O(new_n498));
  nand4 g0113(.a(new_n498), .b(new_n497), .c(new_n496), .d(new_n495), .O(new_n499));
  inv1  g0114(.a(new_n499), .O(new_n500));
  oai21 g0115(.a(\req5 ), .b(new_n495), .c(new_n496), .O(new_n501));
  aoi21 g0116(.a(new_n500), .b(new_n494), .c(new_n501), .O(new_n502));
  inv1  g0117(.a(\priority7 ), .O(new_n503));
  inv1  g0118(.a(\priority8 ), .O(new_n504));
  nor2  g0119(.a(\req8 ), .b(\req7 ), .O(new_n505));
  nand3 g0120(.a(new_n505), .b(new_n504), .c(new_n503), .O(new_n506));
  inv1  g0121(.a(new_n506), .O(new_n507));
  oai21 g0122(.a(new_n502), .b(\req6 ), .c(new_n507), .O(new_n508));
  aoi21 g0123(.a(\req7 ), .b(new_n504), .c(\req8 ), .O(new_n509));
  aoi21 g0124(.a(new_n509), .b(new_n508), .c(\priority9 ), .O(new_n510));
  nor2  g0125(.a(\priority11 ), .b(\priority10 ), .O(new_n511));
  nor2  g0126(.a(\req10 ), .b(\req9 ), .O(new_n512));
  nand2 g0127(.a(new_n512), .b(new_n511), .O(new_n513));
  inv1  g0128(.a(\req10 ), .O(new_n514));
  aoi21 g0129(.a(new_n514), .b(\priority10 ), .c(\priority11 ), .O(new_n515));
  oai21 g0130(.a(new_n513), .b(new_n510), .c(new_n515), .O(new_n516));
  inv1  g0131(.a(\req14 ), .O(new_n517));
  inv1  g0132(.a(\req15 ), .O(new_n518));
  nor2  g0133(.a(\req13 ), .b(\req12 ), .O(new_n519));
  nor2  g0134(.a(\req17 ), .b(\req16 ), .O(new_n520));
  nand4 g0135(.a(new_n520), .b(new_n519), .c(new_n518), .d(new_n517), .O(new_n521));
  nor4  g0136(.a(new_n521), .b(\req18 ), .c(\priority18 ), .d(\priority12 ), .O(new_n522));
  inv1  g0137(.a(new_n522), .O(new_n523));
  aoi21 g0138(.a(new_n516), .b(new_n426), .c(new_n523), .O(new_n524));
  nor2  g0139(.a(\req18 ), .b(\priority18 ), .O(new_n525));
  aoi21 g0140(.a(new_n525), .b(new_n521), .c(\req18 ), .O(new_n526));
  inv1  g0141(.a(new_n526), .O(new_n527));
  oai21 g0142(.a(new_n527), .b(new_n524), .c(new_n425), .O(new_n528));
  inv1  g0143(.a(\priority20 ), .O(new_n529));
  inv1  g0144(.a(\priority21 ), .O(new_n530));
  inv1  g0145(.a(\req19 ), .O(new_n531));
  inv1  g0146(.a(\req20 ), .O(new_n532));
  nand4 g0147(.a(new_n532), .b(new_n531), .c(new_n530), .d(new_n529), .O(new_n533));
  inv1  g0148(.a(new_n533), .O(new_n534));
  aoi21 g0149(.a(new_n532), .b(\priority20 ), .c(\priority21 ), .O(new_n535));
  inv1  g0150(.a(new_n535), .O(new_n536));
  aoi21 g0151(.a(new_n534), .b(new_n528), .c(new_n536), .O(new_n537));
  inv1  g0152(.a(\priority22 ), .O(new_n538));
  inv1  g0153(.a(\priority23 ), .O(new_n539));
  nor2  g0154(.a(\req23 ), .b(\req22 ), .O(new_n540));
  nand3 g0155(.a(new_n540), .b(new_n539), .c(new_n538), .O(new_n541));
  inv1  g0156(.a(new_n541), .O(new_n542));
  oai21 g0157(.a(new_n537), .b(\req21 ), .c(new_n542), .O(new_n543));
  aoi21 g0158(.a(\req22 ), .b(new_n539), .c(\req23 ), .O(new_n544));
  aoi21 g0159(.a(new_n544), .b(new_n543), .c(\priority24 ), .O(new_n545));
  nor2  g0160(.a(\req25 ), .b(\req24 ), .O(new_n546));
  nor2  g0161(.a(\priority26 ), .b(\priority25 ), .O(new_n547));
  nand2 g0162(.a(new_n547), .b(new_n546), .O(new_n548));
  inv1  g0163(.a(\req25 ), .O(new_n549));
  aoi21 g0164(.a(new_n549), .b(\priority25 ), .c(\priority26 ), .O(new_n550));
  oai21 g0165(.a(new_n548), .b(new_n545), .c(new_n550), .O(new_n551));
  inv1  g0166(.a(\priority27 ), .O(new_n552));
  inv1  g0167(.a(\priority28 ), .O(new_n553));
  inv1  g0168(.a(\req27 ), .O(new_n554));
  inv1  g0169(.a(\req28 ), .O(new_n555));
  nand4 g0170(.a(new_n555), .b(new_n554), .c(new_n553), .d(new_n552), .O(new_n556));
  aoi21 g0171(.a(new_n551), .b(new_n424), .c(new_n556), .O(new_n557));
  aoi21 g0172(.a(\req27 ), .b(new_n553), .c(\req28 ), .O(new_n558));
  inv1  g0173(.a(new_n558), .O(new_n559));
  oai21 g0174(.a(new_n559), .b(new_n557), .c(new_n423), .O(new_n560));
  inv1  g0175(.a(\priority30 ), .O(new_n561));
  inv1  g0176(.a(\priority31 ), .O(new_n562));
  inv1  g0177(.a(\req29 ), .O(new_n563));
  inv1  g0178(.a(\req30 ), .O(new_n564));
  nand4 g0179(.a(new_n564), .b(new_n563), .c(new_n562), .d(new_n561), .O(new_n565));
  inv1  g0180(.a(new_n565), .O(new_n566));
  aoi21 g0181(.a(new_n564), .b(\priority30 ), .c(\priority31 ), .O(new_n567));
  inv1  g0182(.a(new_n567), .O(new_n568));
  aoi21 g0183(.a(new_n566), .b(new_n560), .c(new_n568), .O(new_n569));
  inv1  g0184(.a(\req16 ), .O(new_n570));
  aoi21 g0185(.a(new_n570), .b(\priority16 ), .c(\priority17 ), .O(new_n571));
  inv1  g0186(.a(\priority13 ), .O(new_n572));
  nor2  g0187(.a(\priority14 ), .b(new_n572), .O(new_n573));
  nor3  g0188(.a(\req14 ), .b(\req13 ), .c(\priority15 ), .O(new_n574));
  aoi21 g0189(.a(new_n517), .b(\priority14 ), .c(\priority15 ), .O(new_n575));
  inv1  g0190(.a(new_n575), .O(new_n576));
  aoi21 g0191(.a(new_n574), .b(new_n573), .c(new_n576), .O(new_n577));
  nor2  g0192(.a(\req16 ), .b(\priority17 ), .O(new_n578));
  nor2  g0193(.a(\req15 ), .b(\priority16 ), .O(new_n579));
  nand2 g0194(.a(new_n579), .b(new_n578), .O(new_n580));
  oai21 g0195(.a(new_n580), .b(new_n577), .c(new_n571), .O(new_n581));
  inv1  g0196(.a(\req17 ), .O(new_n582));
  inv1  g0197(.a(\req21 ), .O(new_n583));
  nor2  g0198(.a(\req19 ), .b(\req18 ), .O(new_n584));
  nand4 g0199(.a(new_n584), .b(new_n540), .c(new_n583), .d(new_n532), .O(new_n585));
  inv1  g0200(.a(\req31 ), .O(new_n586));
  nand4 g0201(.a(new_n586), .b(new_n564), .c(new_n563), .d(new_n555), .O(new_n587));
  nand3 g0202(.a(new_n546), .b(new_n554), .c(new_n424), .O(new_n588));
  nor3  g0203(.a(new_n588), .b(new_n587), .c(new_n585), .O(new_n589));
  nand2 g0204(.a(new_n589), .b(new_n582), .O(new_n590));
  inv1  g0205(.a(new_n590), .O(new_n591));
  inv1  g0206(.a(\priority32 ), .O(new_n592));
  inv1  g0207(.a(\priority33 ), .O(new_n593));
  inv1  g0208(.a(\req32 ), .O(new_n594));
  inv1  g0209(.a(\req33 ), .O(new_n595));
  nand4 g0210(.a(new_n595), .b(new_n594), .c(new_n593), .d(new_n592), .O(new_n596));
  aoi21 g0211(.a(new_n591), .b(new_n581), .c(new_n596), .O(new_n597));
  oai21 g0212(.a(new_n569), .b(\req31 ), .c(new_n597), .O(new_n598));
  aoi21 g0213(.a(\req32 ), .b(new_n593), .c(\req33 ), .O(new_n599));
  inv1  g0214(.a(\priority34 ), .O(new_n600));
  inv1  g0215(.a(\priority35 ), .O(new_n601));
  inv1  g0216(.a(\req34 ), .O(new_n602));
  inv1  g0217(.a(\req35 ), .O(new_n603));
  nand4 g0218(.a(new_n603), .b(new_n602), .c(new_n601), .d(new_n600), .O(new_n604));
  aoi21 g0219(.a(new_n599), .b(new_n598), .c(new_n604), .O(new_n605));
  aoi21 g0220(.a(\req34 ), .b(new_n601), .c(\req35 ), .O(new_n606));
  inv1  g0221(.a(new_n606), .O(new_n607));
  oai21 g0222(.a(new_n607), .b(new_n605), .c(new_n422), .O(new_n608));
  inv1  g0223(.a(\priority37 ), .O(new_n609));
  inv1  g0224(.a(\priority38 ), .O(new_n610));
  inv1  g0225(.a(\req36 ), .O(new_n611));
  inv1  g0226(.a(\req37 ), .O(new_n612));
  nand4 g0227(.a(new_n612), .b(new_n611), .c(new_n610), .d(new_n609), .O(new_n613));
  inv1  g0228(.a(new_n613), .O(new_n614));
  aoi21 g0229(.a(new_n612), .b(\priority37 ), .c(\priority38 ), .O(new_n615));
  inv1  g0230(.a(new_n615), .O(new_n616));
  aoi21 g0231(.a(new_n614), .b(new_n608), .c(new_n616), .O(new_n617));
  inv1  g0232(.a(\priority39 ), .O(new_n618));
  inv1  g0233(.a(\priority40 ), .O(new_n619));
  inv1  g0234(.a(\req39 ), .O(new_n620));
  inv1  g0235(.a(\req40 ), .O(new_n621));
  nand4 g0236(.a(new_n621), .b(new_n620), .c(new_n619), .d(new_n618), .O(new_n622));
  inv1  g0237(.a(new_n622), .O(new_n623));
  oai21 g0238(.a(new_n617), .b(\req38 ), .c(new_n623), .O(new_n624));
  aoi21 g0239(.a(\req39 ), .b(new_n619), .c(\req40 ), .O(new_n625));
  aoi21 g0240(.a(new_n625), .b(new_n624), .c(\priority41 ), .O(new_n626));
  inv1  g0241(.a(\priority42 ), .O(new_n627));
  inv1  g0242(.a(\priority43 ), .O(new_n628));
  inv1  g0243(.a(\req41 ), .O(new_n629));
  inv1  g0244(.a(\req42 ), .O(new_n630));
  nand4 g0245(.a(new_n630), .b(new_n629), .c(new_n628), .d(new_n627), .O(new_n631));
  aoi21 g0246(.a(new_n630), .b(\priority42 ), .c(\priority43 ), .O(new_n632));
  oai21 g0247(.a(new_n631), .b(new_n626), .c(new_n632), .O(new_n633));
  inv1  g0248(.a(\priority44 ), .O(new_n634));
  inv1  g0249(.a(\priority45 ), .O(new_n635));
  inv1  g0250(.a(\req44 ), .O(new_n636));
  inv1  g0251(.a(\req45 ), .O(new_n637));
  nand4 g0252(.a(new_n637), .b(new_n636), .c(new_n635), .d(new_n634), .O(new_n638));
  aoi21 g0253(.a(new_n633), .b(new_n421), .c(new_n638), .O(new_n639));
  aoi21 g0254(.a(\req44 ), .b(new_n635), .c(\req45 ), .O(new_n640));
  inv1  g0255(.a(new_n640), .O(new_n641));
  oai21 g0256(.a(new_n641), .b(new_n639), .c(new_n420), .O(new_n642));
  inv1  g0257(.a(\priority47 ), .O(new_n643));
  inv1  g0258(.a(\priority48 ), .O(new_n644));
  inv1  g0259(.a(\req46 ), .O(new_n645));
  inv1  g0260(.a(\req47 ), .O(new_n646));
  nand4 g0261(.a(new_n646), .b(new_n645), .c(new_n644), .d(new_n643), .O(new_n647));
  inv1  g0262(.a(new_n647), .O(new_n648));
  aoi21 g0263(.a(new_n646), .b(\priority47 ), .c(\priority48 ), .O(new_n649));
  inv1  g0264(.a(new_n649), .O(new_n650));
  aoi21 g0265(.a(new_n648), .b(new_n642), .c(new_n650), .O(new_n651));
  inv1  g0266(.a(\priority49 ), .O(new_n652));
  inv1  g0267(.a(\priority50 ), .O(new_n653));
  inv1  g0268(.a(\req49 ), .O(new_n654));
  inv1  g0269(.a(\req50 ), .O(new_n655));
  nand4 g0270(.a(new_n655), .b(new_n654), .c(new_n653), .d(new_n652), .O(new_n656));
  inv1  g0271(.a(new_n656), .O(new_n657));
  oai21 g0272(.a(new_n651), .b(\req48 ), .c(new_n657), .O(new_n658));
  aoi21 g0273(.a(\req49 ), .b(new_n653), .c(\req50 ), .O(new_n659));
  aoi21 g0274(.a(new_n659), .b(new_n658), .c(\priority51 ), .O(new_n660));
  inv1  g0275(.a(\priority52 ), .O(new_n661));
  inv1  g0276(.a(\priority53 ), .O(new_n662));
  inv1  g0277(.a(\req51 ), .O(new_n663));
  inv1  g0278(.a(\req52 ), .O(new_n664));
  nand4 g0279(.a(new_n664), .b(new_n663), .c(new_n662), .d(new_n661), .O(new_n665));
  aoi21 g0280(.a(new_n664), .b(\priority52 ), .c(\priority53 ), .O(new_n666));
  oai21 g0281(.a(new_n665), .b(new_n660), .c(new_n666), .O(new_n667));
  inv1  g0282(.a(\priority54 ), .O(new_n668));
  inv1  g0283(.a(\priority55 ), .O(new_n669));
  inv1  g0284(.a(\req54 ), .O(new_n670));
  inv1  g0285(.a(\req55 ), .O(new_n671));
  nand4 g0286(.a(new_n671), .b(new_n670), .c(new_n669), .d(new_n668), .O(new_n672));
  aoi21 g0287(.a(new_n667), .b(new_n419), .c(new_n672), .O(new_n673));
  aoi21 g0288(.a(\req54 ), .b(new_n669), .c(\req55 ), .O(new_n674));
  inv1  g0289(.a(new_n674), .O(new_n675));
  oai21 g0290(.a(new_n675), .b(new_n673), .c(new_n418), .O(new_n676));
  inv1  g0291(.a(\priority57 ), .O(new_n677));
  inv1  g0292(.a(\priority58 ), .O(new_n678));
  inv1  g0293(.a(\req56 ), .O(new_n679));
  inv1  g0294(.a(\req57 ), .O(new_n680));
  nand4 g0295(.a(new_n680), .b(new_n679), .c(new_n678), .d(new_n677), .O(new_n681));
  inv1  g0296(.a(new_n681), .O(new_n682));
  aoi21 g0297(.a(new_n680), .b(\priority57 ), .c(\priority58 ), .O(new_n683));
  inv1  g0298(.a(new_n683), .O(new_n684));
  aoi21 g0299(.a(new_n682), .b(new_n676), .c(new_n684), .O(new_n685));
  inv1  g0300(.a(\priority59 ), .O(new_n686));
  inv1  g0301(.a(\priority60 ), .O(new_n687));
  inv1  g0302(.a(\req59 ), .O(new_n688));
  inv1  g0303(.a(\req60 ), .O(new_n689));
  nand4 g0304(.a(new_n689), .b(new_n688), .c(new_n687), .d(new_n686), .O(new_n690));
  inv1  g0305(.a(new_n690), .O(new_n691));
  oai21 g0306(.a(new_n685), .b(\req58 ), .c(new_n691), .O(new_n692));
  aoi21 g0307(.a(\req59 ), .b(new_n687), .c(\req60 ), .O(new_n693));
  aoi21 g0308(.a(new_n693), .b(new_n692), .c(\priority61 ), .O(new_n694));
  inv1  g0309(.a(\priority73 ), .O(new_n695));
  inv1  g0310(.a(\req72 ), .O(new_n696));
  inv1  g0311(.a(\req69 ), .O(new_n697));
  inv1  g0312(.a(\priority67 ), .O(new_n698));
  aoi21 g0313(.a(new_n406), .b(\priority63 ), .c(\priority64 ), .O(new_n699));
  inv1  g0314(.a(\priority63 ), .O(new_n700));
  inv1  g0315(.a(\req62 ), .O(new_n701));
  nor2  g0316(.a(\req63 ), .b(\priority64 ), .O(new_n702));
  nand4 g0317(.a(new_n702), .b(new_n701), .c(new_n700), .d(\priority62 ), .O(new_n703));
  aoi21 g0318(.a(new_n703), .b(new_n699), .c(\req64 ), .O(new_n704));
  inv1  g0319(.a(\priority65 ), .O(new_n705));
  inv1  g0320(.a(\priority66 ), .O(new_n706));
  nand3 g0321(.a(new_n409), .b(new_n706), .c(new_n705), .O(new_n707));
  aoi21 g0322(.a(\req65 ), .b(new_n706), .c(\req66 ), .O(new_n708));
  oai21 g0323(.a(new_n707), .b(new_n704), .c(new_n708), .O(new_n709));
  inv1  g0324(.a(\priority68 ), .O(new_n710));
  inv1  g0325(.a(\priority69 ), .O(new_n711));
  nand4 g0326(.a(new_n412), .b(new_n411), .c(new_n711), .d(new_n710), .O(new_n712));
  aoi21 g0327(.a(new_n709), .b(new_n698), .c(new_n712), .O(new_n713));
  oai21 g0328(.a(\req68 ), .b(new_n710), .c(new_n711), .O(new_n714));
  oai21 g0329(.a(new_n714), .b(new_n713), .c(new_n697), .O(new_n715));
  inv1  g0330(.a(\priority70 ), .O(new_n716));
  inv1  g0331(.a(\priority71 ), .O(new_n717));
  inv1  g0332(.a(\req70 ), .O(new_n718));
  inv1  g0333(.a(\req71 ), .O(new_n719));
  nand4 g0334(.a(new_n719), .b(new_n718), .c(new_n717), .d(new_n716), .O(new_n720));
  inv1  g0335(.a(new_n720), .O(new_n721));
  oai21 g0336(.a(new_n718), .b(\priority71 ), .c(new_n719), .O(new_n722));
  aoi21 g0337(.a(new_n721), .b(new_n715), .c(new_n722), .O(new_n723));
  oai21 g0338(.a(new_n723), .b(\priority72 ), .c(new_n696), .O(new_n724));
  nor2  g0339(.a(\req73 ), .b(\priority74 ), .O(new_n725));
  inv1  g0340(.a(new_n725), .O(new_n726));
  aoi21 g0341(.a(new_n724), .b(new_n695), .c(new_n726), .O(new_n727));
  oai21 g0342(.a(new_n694), .b(new_n417), .c(new_n727), .O(new_n728));
  inv1  g0343(.a(\priority61 ), .O(new_n729));
  nand2 g0344(.a(new_n693), .b(new_n692), .O(new_n730));
  nand2 g0345(.a(new_n730), .b(new_n729), .O(new_n731));
  aoi21 g0346(.a(new_n731), .b(new_n416), .c(\priority74 ), .O(new_n732));
  aoi21 g0347(.a(new_n732), .b(new_n728), .c(\req74 ), .O(new_n733));
  inv1  g0348(.a(\priority75 ), .O(new_n734));
  inv1  g0349(.a(\priority76 ), .O(new_n735));
  inv1  g0350(.a(\req75 ), .O(new_n736));
  inv1  g0351(.a(\req76 ), .O(new_n737));
  nand4 g0352(.a(new_n737), .b(new_n736), .c(new_n735), .d(new_n734), .O(new_n738));
  aoi21 g0353(.a(\req75 ), .b(new_n735), .c(\req76 ), .O(new_n739));
  oai21 g0354(.a(new_n738), .b(new_n733), .c(new_n739), .O(new_n740));
  inv1  g0355(.a(\priority78 ), .O(new_n741));
  inv1  g0356(.a(\priority79 ), .O(new_n742));
  inv1  g0357(.a(\req77 ), .O(new_n743));
  nand4 g0358(.a(new_n402), .b(new_n743), .c(new_n742), .d(new_n741), .O(new_n744));
  aoi21 g0359(.a(new_n740), .b(new_n405), .c(new_n744), .O(new_n745));
  oai21 g0360(.a(new_n745), .b(new_n404), .c(new_n401), .O(new_n746));
  inv1  g0361(.a(\priority80 ), .O(new_n747));
  inv1  g0362(.a(\priority81 ), .O(new_n748));
  inv1  g0363(.a(\req80 ), .O(new_n749));
  inv1  g0364(.a(\req81 ), .O(new_n750));
  nand4 g0365(.a(new_n750), .b(new_n749), .c(new_n748), .d(new_n747), .O(new_n751));
  inv1  g0366(.a(new_n751), .O(new_n752));
  aoi21 g0367(.a(\req80 ), .b(new_n748), .c(\req81 ), .O(new_n753));
  inv1  g0368(.a(new_n753), .O(new_n754));
  aoi21 g0369(.a(new_n752), .b(new_n746), .c(new_n754), .O(new_n755));
  inv1  g0370(.a(\priority83 ), .O(new_n756));
  inv1  g0371(.a(\priority84 ), .O(new_n757));
  inv1  g0372(.a(\req82 ), .O(new_n758));
  nand4 g0373(.a(new_n399), .b(new_n758), .c(new_n757), .d(new_n756), .O(new_n759));
  inv1  g0374(.a(new_n759), .O(new_n760));
  oai21 g0375(.a(new_n755), .b(\priority82 ), .c(new_n760), .O(new_n761));
  aoi21 g0376(.a(new_n761), .b(new_n400), .c(\req84 ), .O(new_n762));
  inv1  g0377(.a(\priority85 ), .O(new_n763));
  inv1  g0378(.a(\priority86 ), .O(new_n764));
  inv1  g0379(.a(\req85 ), .O(new_n765));
  inv1  g0380(.a(\req86 ), .O(new_n766));
  nand4 g0381(.a(new_n766), .b(new_n765), .c(new_n764), .d(new_n763), .O(new_n767));
  aoi21 g0382(.a(\req85 ), .b(new_n764), .c(\req86 ), .O(new_n768));
  oai21 g0383(.a(new_n767), .b(new_n762), .c(new_n768), .O(new_n769));
  inv1  g0384(.a(\priority88 ), .O(new_n770));
  inv1  g0385(.a(\priority89 ), .O(new_n771));
  inv1  g0386(.a(\req87 ), .O(new_n772));
  nand4 g0387(.a(new_n395), .b(new_n772), .c(new_n771), .d(new_n770), .O(new_n773));
  aoi21 g0388(.a(new_n769), .b(new_n398), .c(new_n773), .O(new_n774));
  oai21 g0389(.a(new_n774), .b(new_n397), .c(new_n394), .O(new_n775));
  inv1  g0390(.a(\priority90 ), .O(new_n776));
  inv1  g0391(.a(\priority91 ), .O(new_n777));
  inv1  g0392(.a(\req90 ), .O(new_n778));
  inv1  g0393(.a(\req91 ), .O(new_n779));
  nand4 g0394(.a(new_n779), .b(new_n778), .c(new_n777), .d(new_n776), .O(new_n780));
  inv1  g0395(.a(new_n780), .O(new_n781));
  aoi21 g0396(.a(\req90 ), .b(new_n777), .c(\req91 ), .O(new_n782));
  inv1  g0397(.a(new_n782), .O(new_n783));
  aoi21 g0398(.a(new_n781), .b(new_n775), .c(new_n783), .O(new_n784));
  nor2  g0399(.a(\req93 ), .b(\priority94 ), .O(new_n785));
  nor2  g0400(.a(\req92 ), .b(\priority93 ), .O(new_n786));
  nand2 g0401(.a(new_n786), .b(new_n785), .O(new_n787));
  inv1  g0402(.a(new_n787), .O(new_n788));
  oai21 g0403(.a(new_n784), .b(\priority92 ), .c(new_n788), .O(new_n789));
  aoi21 g0404(.a(new_n789), .b(new_n393), .c(\req94 ), .O(new_n790));
  inv1  g0405(.a(\priority95 ), .O(new_n791));
  inv1  g0406(.a(\priority96 ), .O(new_n792));
  inv1  g0407(.a(\req95 ), .O(new_n793));
  inv1  g0408(.a(\req96 ), .O(new_n794));
  nand4 g0409(.a(new_n794), .b(new_n793), .c(new_n792), .d(new_n791), .O(new_n795));
  aoi21 g0410(.a(\req95 ), .b(new_n792), .c(\req96 ), .O(new_n796));
  oai21 g0411(.a(new_n795), .b(new_n790), .c(new_n796), .O(new_n797));
  inv1  g0412(.a(\priority98 ), .O(new_n798));
  inv1  g0413(.a(\priority99 ), .O(new_n799));
  nor2  g0414(.a(\req98 ), .b(\req97 ), .O(new_n800));
  nand3 g0415(.a(new_n800), .b(new_n799), .c(new_n798), .O(new_n801));
  aoi21 g0416(.a(new_n797), .b(new_n391), .c(new_n801), .O(new_n802));
  oai21 g0417(.a(\req98 ), .b(new_n798), .c(new_n799), .O(new_n803));
  oai21 g0418(.a(new_n803), .b(new_n802), .c(new_n390), .O(new_n804));
  inv1  g0419(.a(\priority100 ), .O(new_n805));
  inv1  g0420(.a(\priority101 ), .O(new_n806));
  inv1  g0421(.a(\req100 ), .O(new_n807));
  inv1  g0422(.a(\req101 ), .O(new_n808));
  nand4 g0423(.a(new_n808), .b(new_n807), .c(new_n806), .d(new_n805), .O(new_n809));
  inv1  g0424(.a(new_n809), .O(new_n810));
  aoi21 g0425(.a(\req100 ), .b(new_n806), .c(\req101 ), .O(new_n811));
  inv1  g0426(.a(new_n811), .O(new_n812));
  aoi21 g0427(.a(new_n810), .b(new_n804), .c(new_n812), .O(new_n813));
  inv1  g0428(.a(\priority107 ), .O(new_n814));
  inv1  g0429(.a(\priority108 ), .O(new_n815));
  inv1  g0430(.a(\req106 ), .O(new_n816));
  inv1  g0431(.a(\priority104 ), .O(new_n817));
  nor2  g0432(.a(\priority105 ), .b(new_n817), .O(new_n818));
  nor3  g0433(.a(\req105 ), .b(\req104 ), .c(\priority106 ), .O(new_n819));
  nand2 g0434(.a(new_n819), .b(new_n818), .O(new_n820));
  inv1  g0435(.a(\req105 ), .O(new_n821));
  aoi21 g0436(.a(new_n821), .b(\priority105 ), .c(\priority106 ), .O(new_n822));
  nand2 g0437(.a(new_n822), .b(new_n820), .O(new_n823));
  nand2 g0438(.a(new_n823), .b(new_n816), .O(new_n824));
  nor2  g0439(.a(\req108 ), .b(\req107 ), .O(new_n825));
  nand4 g0440(.a(new_n825), .b(new_n824), .c(new_n815), .d(new_n814), .O(new_n826));
  aoi21 g0441(.a(\req107 ), .b(new_n815), .c(\req108 ), .O(new_n827));
  aoi21 g0442(.a(new_n827), .b(new_n826), .c(\priority109 ), .O(new_n828));
  nor2  g0443(.a(\req104 ), .b(\req103 ), .O(new_n829));
  nor2  g0444(.a(\req106 ), .b(\req105 ), .O(new_n830));
  nand3 g0445(.a(new_n830), .b(new_n829), .c(new_n825), .O(new_n831));
  inv1  g0446(.a(new_n831), .O(new_n832));
  nor2  g0447(.a(\req102 ), .b(\priority103 ), .O(new_n833));
  nand3 g0448(.a(new_n833), .b(new_n832), .c(new_n828), .O(new_n834));
  inv1  g0449(.a(new_n834), .O(new_n835));
  oai21 g0450(.a(new_n813), .b(\priority102 ), .c(new_n835), .O(new_n836));
  inv1  g0451(.a(\priority103 ), .O(new_n837));
  oai21 g0452(.a(new_n831), .b(new_n837), .c(new_n828), .O(new_n838));
  inv1  g0453(.a(new_n838), .O(new_n839));
  aoi21 g0454(.a(new_n839), .b(new_n836), .c(\req109 ), .O(new_n840));
  inv1  g0455(.a(\priority110 ), .O(new_n841));
  inv1  g0456(.a(\priority111 ), .O(new_n842));
  inv1  g0457(.a(\req110 ), .O(new_n843));
  inv1  g0458(.a(\req111 ), .O(new_n844));
  nand4 g0459(.a(new_n844), .b(new_n843), .c(new_n842), .d(new_n841), .O(new_n845));
  aoi21 g0460(.a(\req110 ), .b(new_n842), .c(\req111 ), .O(new_n846));
  oai21 g0461(.a(new_n845), .b(new_n840), .c(new_n846), .O(new_n847));
  nor3  g0462(.a(\req113 ), .b(\req112 ), .c(\priority113 ), .O(new_n848));
  nand3 g0463(.a(new_n848), .b(new_n847), .c(new_n389), .O(new_n849));
  aoi21 g0464(.a(\req112 ), .b(new_n449), .c(\req113 ), .O(new_n850));
  nand2 g0465(.a(new_n850), .b(new_n849), .O(new_n851));
  nand2 g0466(.a(new_n851), .b(new_n388), .O(new_n852));
  nor2  g0467(.a(\req114 ), .b(\priority115 ), .O(new_n853));
  nor2  g0468(.a(\req115 ), .b(\priority116 ), .O(new_n854));
  nand3 g0469(.a(new_n854), .b(new_n853), .c(new_n852), .O(new_n855));
  inv1  g0470(.a(\req115 ), .O(new_n856));
  aoi21 g0471(.a(new_n856), .b(\priority115 ), .c(\priority116 ), .O(new_n857));
  nand2 g0472(.a(new_n857), .b(new_n855), .O(new_n858));
  nor2  g0473(.a(\req116 ), .b(\priority117 ), .O(new_n859));
  nor2  g0474(.a(\req117 ), .b(\priority118 ), .O(new_n860));
  nand3 g0475(.a(new_n860), .b(new_n859), .c(new_n858), .O(new_n861));
  aoi21 g0476(.a(new_n435), .b(\priority117 ), .c(\priority118 ), .O(new_n862));
  aoi21 g0477(.a(new_n862), .b(new_n861), .c(\req118 ), .O(new_n863));
  inv1  g0478(.a(\priority120 ), .O(new_n864));
  nand3 g0479(.a(new_n431), .b(new_n864), .c(new_n456), .O(new_n865));
  aoi21 g0480(.a(\req119 ), .b(new_n864), .c(\req120 ), .O(new_n866));
  oai21 g0481(.a(new_n865), .b(new_n863), .c(new_n866), .O(new_n867));
  nand2 g0482(.a(new_n867), .b(new_n387), .O(new_n868));
  inv1  g0483(.a(\priority122 ), .O(new_n869));
  inv1  g0484(.a(\req123 ), .O(new_n870));
  nand4 g0485(.a(new_n870), .b(new_n430), .c(new_n468), .d(new_n869), .O(new_n871));
  inv1  g0486(.a(new_n871), .O(new_n872));
  nand3 g0487(.a(new_n872), .b(new_n868), .c(\req121 ), .O(new_n873));
  nand4 g0488(.a(new_n870), .b(new_n430), .c(new_n468), .d(new_n869), .O(new_n874));
  inv1  g0489(.a(new_n874), .O(new_n875));
  nand3 g0490(.a(new_n875), .b(new_n867), .c(new_n387), .O(new_n876));
  aoi21 g0491(.a(\req122 ), .b(new_n468), .c(\req123 ), .O(new_n877));
  nand3 g0492(.a(new_n877), .b(new_n876), .c(new_n873), .O(new_n878));
  inv1  g0493(.a(\req124 ), .O(new_n879));
  nand4 g0494(.a(new_n475), .b(new_n879), .c(new_n473), .d(new_n469), .O(new_n880));
  inv1  g0495(.a(new_n880), .O(new_n881));
  oai21 g0496(.a(new_n879), .b(\priority125 ), .c(new_n475), .O(new_n882));
  aoi21 g0497(.a(new_n881), .b(new_n878), .c(new_n882), .O(new_n883));
  nor2  g0498(.a(\req126 ), .b(\priority127 ), .O(new_n884));
  oai21 g0499(.a(new_n883), .b(\priority126 ), .c(new_n884), .O(new_n885));
  nor2  g0500(.a(\req127 ), .b(\priority0 ), .O(new_n886));
  inv1  g0501(.a(new_n886), .O(new_n887));
  inv1  g0502(.a(\req127 ), .O(new_n888));
  aoi21 g0503(.a(new_n888), .b(\priority127 ), .c(\priority0 ), .O(new_n889));
  oai21 g0504(.a(new_n887), .b(new_n885), .c(new_n889), .O(new_n890));
  inv1  g0505(.a(new_n890), .O(new_n891));
  nor2  g0506(.a(new_n891), .b(new_n386), .O(\grant0 ));
  inv1  g0507(.a(\priority1 ), .O(new_n893));
  nor2  g0508(.a(new_n891), .b(\req0 ), .O(new_n894));
  inv1  g0509(.a(new_n894), .O(new_n895));
  aoi21 g0510(.a(new_n895), .b(new_n893), .c(new_n428), .O(\grant1 ));
  nand4 g0511(.a(new_n894), .b(new_n428), .c(new_n487), .d(new_n893), .O(new_n897));
  aoi21 g0512(.a(new_n428), .b(\priority1 ), .c(\priority2 ), .O(new_n898));
  aoi21 g0513(.a(new_n898), .b(new_n897), .c(new_n489), .O(\grant2 ));
  nand4 g0514(.a(new_n489), .b(new_n428), .c(new_n487), .d(new_n893), .O(new_n900));
  aoi21 g0515(.a(new_n890), .b(new_n386), .c(new_n900), .O(new_n901));
  aoi21 g0516(.a(\req1 ), .b(new_n487), .c(\req2 ), .O(new_n902));
  inv1  g0517(.a(new_n902), .O(new_n903));
  oai21 g0518(.a(new_n903), .b(new_n901), .c(new_n488), .O(new_n904));
  inv1  g0519(.a(new_n904), .O(new_n905));
  nor2  g0520(.a(new_n905), .b(new_n490), .O(\grant3 ));
  nor2  g0521(.a(\req3 ), .b(\priority4 ), .O(new_n907));
  nand2 g0522(.a(new_n907), .b(new_n904), .O(new_n908));
  aoi21 g0523(.a(new_n908), .b(new_n427), .c(new_n497), .O(\grant4 ));
  nor2  g0524(.a(\req4 ), .b(\priority5 ), .O(new_n910));
  nand3 g0525(.a(new_n910), .b(new_n907), .c(new_n904), .O(new_n911));
  aoi21 g0526(.a(new_n497), .b(\priority4 ), .c(\priority5 ), .O(new_n912));
  aoi21 g0527(.a(new_n912), .b(new_n911), .c(new_n498), .O(\grant5 ));
  inv1  g0528(.a(\req6 ), .O(new_n914));
  aoi21 g0529(.a(new_n912), .b(new_n911), .c(\req5 ), .O(new_n915));
  inv1  g0530(.a(new_n915), .O(new_n916));
  aoi21 g0531(.a(new_n916), .b(new_n496), .c(new_n914), .O(\grant6 ));
  inv1  g0532(.a(\req7 ), .O(new_n918));
  nand4 g0533(.a(new_n915), .b(new_n914), .c(new_n503), .d(new_n496), .O(new_n919));
  aoi21 g0534(.a(new_n914), .b(\priority6 ), .c(\priority7 ), .O(new_n920));
  aoi21 g0535(.a(new_n920), .b(new_n919), .c(new_n918), .O(\grant7 ));
  inv1  g0536(.a(\req8 ), .O(new_n922));
  nand4 g0537(.a(new_n918), .b(new_n914), .c(new_n503), .d(new_n496), .O(new_n923));
  aoi21 g0538(.a(\req6 ), .b(new_n503), .c(\req7 ), .O(new_n924));
  oai21 g0539(.a(new_n923), .b(new_n915), .c(new_n924), .O(new_n925));
  aoi21 g0540(.a(new_n925), .b(new_n504), .c(new_n922), .O(\grant8 ));
  inv1  g0541(.a(\req9 ), .O(new_n927));
  nand2 g0542(.a(new_n925), .b(new_n504), .O(new_n928));
  aoi21 g0543(.a(new_n928), .b(new_n922), .c(\priority9 ), .O(new_n929));
  nor2  g0544(.a(new_n929), .b(new_n927), .O(\grant9 ));
  nor2  g0545(.a(\req8 ), .b(\priority9 ), .O(new_n931));
  nor2  g0546(.a(\req9 ), .b(\priority10 ), .O(new_n932));
  nand3 g0547(.a(new_n932), .b(new_n931), .c(new_n928), .O(new_n933));
  aoi21 g0548(.a(new_n927), .b(\priority9 ), .c(\priority10 ), .O(new_n934));
  aoi21 g0549(.a(new_n934), .b(new_n933), .c(new_n514), .O(\grant10 ));
  nand2 g0550(.a(new_n934), .b(new_n933), .O(new_n936));
  aoi21 g0551(.a(new_n936), .b(new_n514), .c(\priority11 ), .O(new_n937));
  nor2  g0552(.a(new_n937), .b(new_n426), .O(\grant11 ));
  inv1  g0553(.a(\req12 ), .O(new_n939));
  nor2  g0554(.a(\req10 ), .b(\priority11 ), .O(new_n940));
  nor2  g0555(.a(\req11 ), .b(\priority12 ), .O(new_n941));
  nand3 g0556(.a(new_n941), .b(new_n940), .c(new_n936), .O(new_n942));
  aoi21 g0557(.a(new_n426), .b(\priority11 ), .c(\priority12 ), .O(new_n943));
  aoi21 g0558(.a(new_n943), .b(new_n942), .c(new_n939), .O(\grant12 ));
  inv1  g0559(.a(\req13 ), .O(new_n945));
  aoi21 g0560(.a(new_n943), .b(new_n942), .c(\req12 ), .O(new_n946));
  inv1  g0561(.a(new_n946), .O(new_n947));
  aoi21 g0562(.a(new_n947), .b(new_n572), .c(new_n945), .O(\grant13 ));
  inv1  g0563(.a(\priority14 ), .O(new_n949));
  nand4 g0564(.a(new_n946), .b(new_n945), .c(new_n949), .d(new_n572), .O(new_n950));
  aoi21 g0565(.a(new_n945), .b(\priority13 ), .c(\priority14 ), .O(new_n951));
  aoi21 g0566(.a(new_n951), .b(new_n950), .c(new_n517), .O(\grant14 ));
  inv1  g0567(.a(\priority15 ), .O(new_n953));
  nand4 g0568(.a(new_n517), .b(new_n945), .c(new_n949), .d(new_n572), .O(new_n954));
  aoi21 g0569(.a(\req13 ), .b(new_n949), .c(\req14 ), .O(new_n955));
  oai21 g0570(.a(new_n954), .b(new_n946), .c(new_n955), .O(new_n956));
  aoi21 g0571(.a(new_n956), .b(new_n953), .c(new_n518), .O(\grant15 ));
  inv1  g0572(.a(\priority16 ), .O(new_n958));
  nand2 g0573(.a(new_n956), .b(new_n953), .O(new_n959));
  nand2 g0574(.a(new_n959), .b(new_n579), .O(new_n960));
  aoi21 g0575(.a(new_n960), .b(new_n958), .c(new_n570), .O(\grant16 ));
  nand3 g0576(.a(new_n959), .b(new_n579), .c(new_n578), .O(new_n962));
  aoi21 g0577(.a(new_n962), .b(new_n571), .c(new_n582), .O(\grant17 ));
  inv1  g0578(.a(\req18 ), .O(new_n964));
  inv1  g0579(.a(\priority17 ), .O(new_n965));
  nand2 g0580(.a(new_n579), .b(new_n570), .O(new_n966));
  aoi21 g0581(.a(\req15 ), .b(new_n958), .c(\req16 ), .O(new_n967));
  oai21 g0582(.a(new_n966), .b(new_n959), .c(new_n967), .O(new_n968));
  nand2 g0583(.a(new_n968), .b(new_n965), .O(new_n969));
  aoi21 g0584(.a(new_n969), .b(new_n582), .c(\priority18 ), .O(new_n970));
  nor2  g0585(.a(new_n970), .b(new_n964), .O(\grant18 ));
  aoi21 g0586(.a(new_n962), .b(new_n571), .c(\req17 ), .O(new_n972));
  nand3 g0587(.a(new_n972), .b(new_n525), .c(new_n425), .O(new_n973));
  aoi21 g0588(.a(new_n964), .b(\priority18 ), .c(\priority19 ), .O(new_n974));
  aoi21 g0589(.a(new_n974), .b(new_n973), .c(new_n531), .O(\grant19 ));
  nand3 g0590(.a(new_n525), .b(new_n531), .c(new_n425), .O(new_n976));
  aoi21 g0591(.a(\req18 ), .b(new_n425), .c(\req19 ), .O(new_n977));
  oai21 g0592(.a(new_n976), .b(new_n972), .c(new_n977), .O(new_n978));
  aoi21 g0593(.a(new_n978), .b(new_n529), .c(new_n532), .O(\grant20 ));
  nand2 g0594(.a(new_n978), .b(new_n529), .O(new_n980));
  aoi21 g0595(.a(new_n980), .b(new_n532), .c(\priority21 ), .O(new_n981));
  nor2  g0596(.a(new_n981), .b(new_n583), .O(\grant21 ));
  inv1  g0597(.a(\req22 ), .O(new_n983));
  nor2  g0598(.a(\req21 ), .b(\priority22 ), .O(new_n984));
  nand4 g0599(.a(new_n984), .b(new_n980), .c(new_n532), .d(new_n530), .O(new_n985));
  aoi21 g0600(.a(new_n583), .b(\priority21 ), .c(\priority22 ), .O(new_n986));
  aoi21 g0601(.a(new_n986), .b(new_n985), .c(new_n983), .O(\grant22 ));
  inv1  g0602(.a(\req23 ), .O(new_n988));
  nand3 g0603(.a(new_n984), .b(new_n983), .c(new_n530), .O(new_n989));
  inv1  g0604(.a(new_n989), .O(new_n990));
  nand3 g0605(.a(new_n990), .b(new_n980), .c(\req20 ), .O(new_n991));
  nand4 g0606(.a(new_n983), .b(new_n583), .c(new_n538), .d(new_n530), .O(new_n992));
  inv1  g0607(.a(new_n992), .O(new_n993));
  nand3 g0608(.a(new_n993), .b(new_n978), .c(new_n529), .O(new_n994));
  aoi21 g0609(.a(\req21 ), .b(new_n538), .c(\req22 ), .O(new_n995));
  nand3 g0610(.a(new_n995), .b(new_n994), .c(new_n991), .O(new_n996));
  aoi21 g0611(.a(new_n996), .b(new_n539), .c(new_n988), .O(\grant23 ));
  inv1  g0612(.a(\req24 ), .O(new_n998));
  inv1  g0613(.a(\priority24 ), .O(new_n999));
  inv1  g0614(.a(new_n996), .O(new_n1000));
  nand4 g0615(.a(new_n1000), .b(new_n988), .c(new_n999), .d(new_n539), .O(new_n1001));
  aoi21 g0616(.a(new_n988), .b(\priority23 ), .c(\priority24 ), .O(new_n1002));
  aoi21 g0617(.a(new_n1002), .b(new_n1001), .c(new_n998), .O(\grant24 ));
  nand4 g0618(.a(new_n998), .b(new_n988), .c(new_n999), .d(new_n539), .O(new_n1004));
  inv1  g0619(.a(new_n1004), .O(new_n1005));
  oai21 g0620(.a(new_n988), .b(\priority24 ), .c(new_n998), .O(new_n1006));
  aoi21 g0621(.a(new_n1005), .b(new_n996), .c(new_n1006), .O(new_n1007));
  nor2  g0622(.a(new_n1007), .b(\priority25 ), .O(new_n1008));
  nor2  g0623(.a(new_n1008), .b(new_n549), .O(\grant25 ));
  inv1  g0624(.a(\priority26 ), .O(new_n1010));
  nor2  g0625(.a(\req25 ), .b(\priority26 ), .O(new_n1011));
  oai21 g0626(.a(new_n1007), .b(\priority25 ), .c(new_n1011), .O(new_n1012));
  aoi21 g0627(.a(new_n1012), .b(new_n1010), .c(new_n424), .O(\grant26 ));
  nor2  g0628(.a(\req26 ), .b(\priority27 ), .O(new_n1014));
  inv1  g0629(.a(new_n1014), .O(new_n1015));
  aoi21 g0630(.a(new_n424), .b(\priority26 ), .c(\priority27 ), .O(new_n1016));
  oai21 g0631(.a(new_n1015), .b(new_n1012), .c(new_n1016), .O(new_n1017));
  inv1  g0632(.a(new_n1017), .O(new_n1018));
  nor2  g0633(.a(new_n1018), .b(new_n554), .O(\grant27 ));
  nand2 g0634(.a(new_n1017), .b(new_n554), .O(new_n1020));
  aoi21 g0635(.a(new_n1020), .b(new_n553), .c(new_n555), .O(\grant28 ));
  nor2  g0636(.a(\req28 ), .b(\priority29 ), .O(new_n1022));
  nand4 g0637(.a(new_n1022), .b(new_n1017), .c(new_n554), .d(new_n553), .O(new_n1023));
  aoi21 g0638(.a(new_n555), .b(\priority28 ), .c(\priority29 ), .O(new_n1024));
  aoi21 g0639(.a(new_n1024), .b(new_n1023), .c(new_n563), .O(\grant29 ));
  nand4 g0640(.a(new_n563), .b(new_n555), .c(new_n423), .d(new_n553), .O(new_n1026));
  aoi21 g0641(.a(new_n1017), .b(new_n554), .c(new_n1026), .O(new_n1027));
  aoi21 g0642(.a(\req28 ), .b(new_n423), .c(\req29 ), .O(new_n1028));
  inv1  g0643(.a(new_n1028), .O(new_n1029));
  oai21 g0644(.a(new_n1029), .b(new_n1027), .c(new_n561), .O(new_n1030));
  inv1  g0645(.a(new_n1030), .O(new_n1031));
  nor2  g0646(.a(new_n1031), .b(new_n564), .O(\grant30 ));
  nor3  g0647(.a(new_n1031), .b(\req30 ), .c(\priority31 ), .O(new_n1033));
  inv1  g0648(.a(new_n1033), .O(new_n1034));
  aoi21 g0649(.a(new_n1034), .b(new_n562), .c(new_n586), .O(\grant31 ));
  nand3 g0650(.a(new_n1033), .b(new_n586), .c(new_n592), .O(new_n1036));
  aoi21 g0651(.a(new_n586), .b(\priority31 ), .c(\priority32 ), .O(new_n1037));
  aoi21 g0652(.a(new_n1037), .b(new_n1036), .c(new_n594), .O(\grant32 ));
  nand4 g0653(.a(new_n594), .b(new_n586), .c(new_n592), .d(new_n562), .O(new_n1039));
  inv1  g0654(.a(new_n1039), .O(new_n1040));
  nand3 g0655(.a(new_n1040), .b(new_n1030), .c(\req30 ), .O(new_n1041));
  inv1  g0656(.a(new_n1026), .O(new_n1042));
  nand2 g0657(.a(new_n1042), .b(new_n1020), .O(new_n1043));
  nand2 g0658(.a(new_n1028), .b(new_n1043), .O(new_n1044));
  nand4 g0659(.a(new_n594), .b(new_n586), .c(new_n592), .d(new_n562), .O(new_n1045));
  inv1  g0660(.a(new_n1045), .O(new_n1046));
  nand3 g0661(.a(new_n1046), .b(new_n1044), .c(new_n561), .O(new_n1047));
  aoi21 g0662(.a(\req31 ), .b(new_n592), .c(\req32 ), .O(new_n1048));
  nand3 g0663(.a(new_n1048), .b(new_n1047), .c(new_n1041), .O(new_n1049));
  aoi21 g0664(.a(new_n1049), .b(new_n593), .c(new_n595), .O(\grant33 ));
  inv1  g0665(.a(new_n1049), .O(new_n1051));
  nand4 g0666(.a(new_n1051), .b(new_n595), .c(new_n600), .d(new_n593), .O(new_n1052));
  aoi21 g0667(.a(new_n595), .b(\priority33 ), .c(\priority34 ), .O(new_n1053));
  aoi21 g0668(.a(new_n1053), .b(new_n1052), .c(new_n602), .O(\grant34 ));
  nand3 g0669(.a(new_n602), .b(new_n595), .c(new_n601), .O(new_n1055));
  nor3  g0670(.a(new_n1055), .b(\priority34 ), .c(new_n593), .O(new_n1056));
  nand2 g0671(.a(new_n1056), .b(new_n1049), .O(new_n1057));
  nand4 g0672(.a(new_n602), .b(new_n595), .c(new_n601), .d(new_n600), .O(new_n1058));
  inv1  g0673(.a(new_n1058), .O(new_n1059));
  nand4 g0674(.a(new_n1059), .b(new_n1048), .c(new_n1047), .d(new_n1041), .O(new_n1060));
  aoi21 g0675(.a(new_n602), .b(\priority34 ), .c(\priority35 ), .O(new_n1061));
  nand3 g0676(.a(new_n1061), .b(new_n1060), .c(new_n1057), .O(new_n1062));
  inv1  g0677(.a(new_n1062), .O(new_n1063));
  nor2  g0678(.a(new_n1063), .b(new_n603), .O(\grant35 ));
  nor3  g0679(.a(new_n1063), .b(\req35 ), .c(\priority36 ), .O(new_n1065));
  inv1  g0680(.a(new_n1065), .O(new_n1066));
  aoi21 g0681(.a(new_n1066), .b(new_n422), .c(new_n611), .O(\grant36 ));
  nand3 g0682(.a(new_n1065), .b(new_n611), .c(new_n609), .O(new_n1068));
  aoi21 g0683(.a(new_n611), .b(\priority36 ), .c(\priority37 ), .O(new_n1069));
  aoi21 g0684(.a(new_n1069), .b(new_n1068), .c(new_n612), .O(\grant37 ));
  inv1  g0685(.a(\req38 ), .O(new_n1071));
  nand4 g0686(.a(new_n612), .b(new_n611), .c(new_n609), .d(new_n422), .O(new_n1072));
  inv1  g0687(.a(new_n1072), .O(new_n1073));
  nand3 g0688(.a(new_n1073), .b(new_n1062), .c(\req35 ), .O(new_n1074));
  nand4 g0689(.a(new_n612), .b(new_n611), .c(new_n609), .d(new_n422), .O(new_n1075));
  inv1  g0690(.a(new_n1075), .O(new_n1076));
  nand4 g0691(.a(new_n1076), .b(new_n1061), .c(new_n1060), .d(new_n1057), .O(new_n1077));
  aoi21 g0692(.a(\req36 ), .b(new_n609), .c(\req37 ), .O(new_n1078));
  nand3 g0693(.a(new_n1078), .b(new_n1077), .c(new_n1074), .O(new_n1079));
  aoi21 g0694(.a(new_n1079), .b(new_n610), .c(new_n1071), .O(\grant38 ));
  inv1  g0695(.a(new_n1079), .O(new_n1081));
  nand4 g0696(.a(new_n1081), .b(new_n1071), .c(new_n618), .d(new_n610), .O(new_n1082));
  aoi21 g0697(.a(new_n1071), .b(\priority38 ), .c(\priority39 ), .O(new_n1083));
  aoi21 g0698(.a(new_n1083), .b(new_n1082), .c(new_n620), .O(\grant39 ));
  nand4 g0699(.a(new_n620), .b(new_n1071), .c(new_n618), .d(new_n610), .O(new_n1085));
  inv1  g0700(.a(new_n1085), .O(new_n1086));
  aoi21 g0701(.a(\req38 ), .b(new_n618), .c(\req39 ), .O(new_n1087));
  inv1  g0702(.a(new_n1087), .O(new_n1088));
  aoi21 g0703(.a(new_n1086), .b(new_n1079), .c(new_n1088), .O(new_n1089));
  nor2  g0704(.a(new_n1089), .b(\priority40 ), .O(new_n1090));
  nor2  g0705(.a(new_n1090), .b(new_n621), .O(\grant40 ));
  inv1  g0706(.a(\priority41 ), .O(new_n1092));
  nor2  g0707(.a(\req40 ), .b(\priority41 ), .O(new_n1093));
  oai21 g0708(.a(new_n1089), .b(\priority40 ), .c(new_n1093), .O(new_n1094));
  aoi21 g0709(.a(new_n1094), .b(new_n1092), .c(new_n629), .O(\grant41 ));
  nor2  g0710(.a(\req41 ), .b(\priority42 ), .O(new_n1096));
  inv1  g0711(.a(new_n1096), .O(new_n1097));
  aoi21 g0712(.a(new_n629), .b(\priority41 ), .c(\priority42 ), .O(new_n1098));
  oai21 g0713(.a(new_n1097), .b(new_n1094), .c(new_n1098), .O(new_n1099));
  inv1  g0714(.a(new_n1099), .O(new_n1100));
  nor2  g0715(.a(new_n1100), .b(new_n630), .O(\grant42 ));
  nor2  g0716(.a(new_n1100), .b(\req42 ), .O(new_n1102));
  inv1  g0717(.a(new_n1102), .O(new_n1103));
  aoi21 g0718(.a(new_n1103), .b(new_n628), .c(new_n421), .O(\grant43 ));
  nand4 g0719(.a(new_n1102), .b(new_n421), .c(new_n634), .d(new_n628), .O(new_n1105));
  aoi21 g0720(.a(new_n421), .b(\priority43 ), .c(\priority44 ), .O(new_n1106));
  aoi21 g0721(.a(new_n1106), .b(new_n1105), .c(new_n636), .O(\grant44 ));
  nand4 g0722(.a(new_n636), .b(new_n421), .c(new_n634), .d(new_n628), .O(new_n1108));
  aoi21 g0723(.a(new_n1099), .b(new_n630), .c(new_n1108), .O(new_n1109));
  aoi21 g0724(.a(\req43 ), .b(new_n634), .c(\req44 ), .O(new_n1110));
  inv1  g0725(.a(new_n1110), .O(new_n1111));
  oai21 g0726(.a(new_n1111), .b(new_n1109), .c(new_n635), .O(new_n1112));
  inv1  g0727(.a(new_n1112), .O(new_n1113));
  nor2  g0728(.a(new_n1113), .b(new_n637), .O(\grant45 ));
  nor2  g0729(.a(\req45 ), .b(\priority46 ), .O(new_n1115));
  nand2 g0730(.a(new_n1115), .b(new_n1112), .O(new_n1116));
  aoi21 g0731(.a(new_n1116), .b(new_n420), .c(new_n645), .O(\grant46 ));
  nor2  g0732(.a(\req46 ), .b(\priority47 ), .O(new_n1118));
  nand3 g0733(.a(new_n1118), .b(new_n1115), .c(new_n1112), .O(new_n1119));
  aoi21 g0734(.a(new_n645), .b(\priority46 ), .c(\priority47 ), .O(new_n1120));
  aoi21 g0735(.a(new_n1120), .b(new_n1119), .c(new_n646), .O(\grant47 ));
  inv1  g0736(.a(\req48 ), .O(new_n1122));
  aoi21 g0737(.a(new_n1120), .b(new_n1119), .c(\req47 ), .O(new_n1123));
  inv1  g0738(.a(new_n1123), .O(new_n1124));
  aoi21 g0739(.a(new_n1124), .b(new_n644), .c(new_n1122), .O(\grant48 ));
  nand4 g0740(.a(new_n1123), .b(new_n1122), .c(new_n652), .d(new_n644), .O(new_n1126));
  aoi21 g0741(.a(new_n1122), .b(\priority48 ), .c(\priority49 ), .O(new_n1127));
  aoi21 g0742(.a(new_n1127), .b(new_n1126), .c(new_n654), .O(\grant49 ));
  nand4 g0743(.a(new_n654), .b(new_n1122), .c(new_n652), .d(new_n644), .O(new_n1129));
  aoi21 g0744(.a(\req48 ), .b(new_n652), .c(\req49 ), .O(new_n1130));
  oai21 g0745(.a(new_n1129), .b(new_n1123), .c(new_n1130), .O(new_n1131));
  aoi21 g0746(.a(new_n1131), .b(new_n653), .c(new_n655), .O(\grant50 ));
  nand2 g0747(.a(new_n1131), .b(new_n653), .O(new_n1133));
  aoi21 g0748(.a(new_n1133), .b(new_n655), .c(\priority51 ), .O(new_n1134));
  nor2  g0749(.a(new_n1134), .b(new_n663), .O(\grant51 ));
  nor2  g0750(.a(\req50 ), .b(\priority51 ), .O(new_n1136));
  nor2  g0751(.a(\req51 ), .b(\priority52 ), .O(new_n1137));
  nand3 g0752(.a(new_n1137), .b(new_n1136), .c(new_n1133), .O(new_n1138));
  aoi21 g0753(.a(new_n663), .b(\priority51 ), .c(\priority52 ), .O(new_n1139));
  aoi21 g0754(.a(new_n1139), .b(new_n1138), .c(new_n664), .O(\grant52 ));
  aoi21 g0755(.a(new_n1139), .b(new_n1138), .c(\req52 ), .O(new_n1141));
  inv1  g0756(.a(new_n1141), .O(new_n1142));
  aoi21 g0757(.a(new_n1142), .b(new_n662), .c(new_n419), .O(\grant53 ));
  nand4 g0758(.a(new_n1141), .b(new_n419), .c(new_n668), .d(new_n662), .O(new_n1144));
  aoi21 g0759(.a(new_n419), .b(\priority53 ), .c(\priority54 ), .O(new_n1145));
  aoi21 g0760(.a(new_n1145), .b(new_n1144), .c(new_n670), .O(\grant54 ));
  nor2  g0761(.a(\req54 ), .b(\req53 ), .O(new_n1147));
  nand3 g0762(.a(new_n1147), .b(new_n668), .c(new_n662), .O(new_n1148));
  aoi21 g0763(.a(\req53 ), .b(new_n668), .c(\req54 ), .O(new_n1149));
  oai21 g0764(.a(new_n1148), .b(new_n1141), .c(new_n1149), .O(new_n1150));
  aoi21 g0765(.a(new_n1150), .b(new_n669), .c(new_n671), .O(\grant55 ));
  nand2 g0766(.a(new_n1150), .b(new_n669), .O(new_n1152));
  nor2  g0767(.a(\req55 ), .b(\priority56 ), .O(new_n1153));
  nand2 g0768(.a(new_n1153), .b(new_n1152), .O(new_n1154));
  aoi21 g0769(.a(new_n1154), .b(new_n418), .c(new_n679), .O(\grant56 ));
  nor2  g0770(.a(\req56 ), .b(\priority57 ), .O(new_n1156));
  nand3 g0771(.a(new_n1156), .b(new_n1153), .c(new_n1152), .O(new_n1157));
  aoi21 g0772(.a(new_n679), .b(\priority56 ), .c(\priority57 ), .O(new_n1158));
  aoi21 g0773(.a(new_n1158), .b(new_n1157), .c(new_n680), .O(\grant57 ));
  inv1  g0774(.a(\req58 ), .O(new_n1160));
  aoi21 g0775(.a(new_n1158), .b(new_n1157), .c(\req57 ), .O(new_n1161));
  inv1  g0776(.a(new_n1161), .O(new_n1162));
  aoi21 g0777(.a(new_n1162), .b(new_n678), .c(new_n1160), .O(\grant58 ));
  nand4 g0778(.a(new_n1161), .b(new_n1160), .c(new_n686), .d(new_n678), .O(new_n1164));
  aoi21 g0779(.a(new_n1160), .b(\priority58 ), .c(\priority59 ), .O(new_n1165));
  aoi21 g0780(.a(new_n1165), .b(new_n1164), .c(new_n688), .O(\grant59 ));
  nand4 g0781(.a(new_n688), .b(new_n1160), .c(new_n686), .d(new_n678), .O(new_n1167));
  aoi21 g0782(.a(\req58 ), .b(new_n686), .c(\req59 ), .O(new_n1168));
  oai21 g0783(.a(new_n1167), .b(new_n1161), .c(new_n1168), .O(new_n1169));
  aoi21 g0784(.a(new_n1169), .b(new_n687), .c(new_n689), .O(\grant60 ));
  inv1  g0785(.a(\req61 ), .O(new_n1171));
  nand2 g0786(.a(new_n1169), .b(new_n687), .O(new_n1172));
  nor2  g0787(.a(\req60 ), .b(\priority61 ), .O(new_n1173));
  nand2 g0788(.a(new_n1173), .b(new_n1172), .O(new_n1174));
  aoi21 g0789(.a(new_n1174), .b(new_n729), .c(new_n1171), .O(\grant61 ));
  inv1  g0790(.a(\priority62 ), .O(new_n1176));
  nand4 g0791(.a(new_n1173), .b(new_n1172), .c(new_n1171), .d(new_n1176), .O(new_n1177));
  aoi21 g0792(.a(new_n1171), .b(\priority61 ), .c(\priority62 ), .O(new_n1178));
  aoi21 g0793(.a(new_n1178), .b(new_n1177), .c(new_n701), .O(\grant62 ));
  nor3  g0794(.a(\req61 ), .b(\req60 ), .c(\priority61 ), .O(new_n1180));
  nand3 g0795(.a(new_n1180), .b(new_n1169), .c(new_n687), .O(new_n1181));
  aoi21 g0796(.a(\req60 ), .b(new_n729), .c(\req61 ), .O(new_n1182));
  nand2 g0797(.a(new_n1182), .b(new_n1181), .O(new_n1183));
  nand2 g0798(.a(new_n1183), .b(new_n1176), .O(new_n1184));
  nor2  g0799(.a(\req62 ), .b(\priority63 ), .O(new_n1185));
  nand2 g0800(.a(new_n1185), .b(new_n1184), .O(new_n1186));
  aoi21 g0801(.a(new_n1186), .b(new_n700), .c(new_n406), .O(\grant63 ));
  nand3 g0802(.a(new_n1185), .b(new_n1184), .c(new_n702), .O(new_n1188));
  aoi21 g0803(.a(new_n1188), .b(new_n699), .c(new_n407), .O(\grant64 ));
  inv1  g0804(.a(\req65 ), .O(new_n1190));
  nand2 g0805(.a(new_n1188), .b(new_n699), .O(new_n1191));
  nor2  g0806(.a(\req64 ), .b(\priority65 ), .O(new_n1192));
  nand2 g0807(.a(new_n1192), .b(new_n1191), .O(new_n1193));
  aoi21 g0808(.a(new_n1193), .b(new_n705), .c(new_n1190), .O(\grant65 ));
  inv1  g0809(.a(\req66 ), .O(new_n1195));
  nor2  g0810(.a(\req65 ), .b(\priority66 ), .O(new_n1196));
  nand3 g0811(.a(new_n1196), .b(new_n1192), .c(new_n1191), .O(new_n1197));
  aoi21 g0812(.a(new_n1190), .b(\priority65 ), .c(\priority66 ), .O(new_n1198));
  aoi21 g0813(.a(new_n1198), .b(new_n1197), .c(new_n1195), .O(\grant66 ));
  nand2 g0814(.a(new_n1198), .b(new_n1197), .O(new_n1200));
  nor2  g0815(.a(\req66 ), .b(\priority67 ), .O(new_n1201));
  nand2 g0816(.a(new_n1201), .b(new_n1200), .O(new_n1202));
  aoi21 g0817(.a(new_n1202), .b(new_n698), .c(new_n411), .O(\grant67 ));
  nor2  g0818(.a(\req67 ), .b(\priority68 ), .O(new_n1204));
  nand3 g0819(.a(new_n1204), .b(new_n1201), .c(new_n1200), .O(new_n1205));
  aoi21 g0820(.a(new_n411), .b(\priority67 ), .c(\priority68 ), .O(new_n1206));
  aoi21 g0821(.a(new_n1206), .b(new_n1205), .c(new_n412), .O(\grant68 ));
  nand2 g0822(.a(new_n1206), .b(new_n1205), .O(new_n1208));
  nor2  g0823(.a(\req68 ), .b(\priority69 ), .O(new_n1209));
  nand2 g0824(.a(new_n1209), .b(new_n1208), .O(new_n1210));
  aoi21 g0825(.a(new_n1210), .b(new_n711), .c(new_n697), .O(\grant69 ));
  nor2  g0826(.a(\req69 ), .b(\priority70 ), .O(new_n1212));
  nand3 g0827(.a(new_n1212), .b(new_n1209), .c(new_n1208), .O(new_n1213));
  aoi21 g0828(.a(new_n697), .b(\priority69 ), .c(\priority70 ), .O(new_n1214));
  aoi21 g0829(.a(new_n1214), .b(new_n1213), .c(new_n718), .O(\grant70 ));
  nand2 g0830(.a(new_n1214), .b(new_n1213), .O(new_n1216));
  nor2  g0831(.a(\req70 ), .b(\priority71 ), .O(new_n1217));
  nand2 g0832(.a(new_n1217), .b(new_n1216), .O(new_n1218));
  aoi21 g0833(.a(new_n1218), .b(new_n717), .c(new_n719), .O(\grant71 ));
  nor2  g0834(.a(\req71 ), .b(\priority72 ), .O(new_n1220));
  nand3 g0835(.a(new_n1220), .b(new_n1217), .c(new_n1216), .O(new_n1221));
  aoi21 g0836(.a(new_n719), .b(\priority71 ), .c(\priority72 ), .O(new_n1222));
  aoi21 g0837(.a(new_n1222), .b(new_n1221), .c(new_n696), .O(\grant72 ));
  inv1  g0838(.a(\req73 ), .O(new_n1224));
  aoi21 g0839(.a(new_n1222), .b(new_n1221), .c(\req72 ), .O(new_n1225));
  inv1  g0840(.a(new_n1225), .O(new_n1226));
  aoi21 g0841(.a(new_n1226), .b(new_n695), .c(new_n1224), .O(\grant73 ));
  inv1  g0842(.a(\req74 ), .O(new_n1228));
  nand3 g0843(.a(new_n1225), .b(new_n725), .c(new_n695), .O(new_n1229));
  aoi21 g0844(.a(new_n1224), .b(\priority73 ), .c(\priority74 ), .O(new_n1230));
  aoi21 g0845(.a(new_n1230), .b(new_n1229), .c(new_n1228), .O(\grant74 ));
  inv1  g0846(.a(\priority74 ), .O(new_n1232));
  nand4 g0847(.a(new_n1228), .b(new_n1224), .c(new_n1232), .d(new_n695), .O(new_n1233));
  aoi21 g0848(.a(\req73 ), .b(new_n1232), .c(\req74 ), .O(new_n1234));
  oai21 g0849(.a(new_n1233), .b(new_n1225), .c(new_n1234), .O(new_n1235));
  aoi21 g0850(.a(new_n1235), .b(new_n734), .c(new_n736), .O(\grant75 ));
  nand2 g0851(.a(new_n1235), .b(new_n734), .O(new_n1237));
  nor2  g0852(.a(\req75 ), .b(\priority76 ), .O(new_n1238));
  nand2 g0853(.a(new_n1238), .b(new_n1237), .O(new_n1239));
  aoi21 g0854(.a(new_n1239), .b(new_n735), .c(new_n737), .O(\grant76 ));
  nor2  g0855(.a(\req76 ), .b(\priority77 ), .O(new_n1241));
  nand3 g0856(.a(new_n1241), .b(new_n1238), .c(new_n1237), .O(new_n1242));
  aoi21 g0857(.a(new_n737), .b(\priority76 ), .c(\priority77 ), .O(new_n1243));
  aoi21 g0858(.a(new_n1243), .b(new_n1242), .c(new_n743), .O(\grant77 ));
  aoi21 g0859(.a(new_n1243), .b(new_n1242), .c(\req77 ), .O(new_n1245));
  inv1  g0860(.a(new_n1245), .O(new_n1246));
  aoi21 g0861(.a(new_n1246), .b(new_n741), .c(new_n402), .O(\grant78 ));
  nand4 g0862(.a(new_n1245), .b(new_n402), .c(new_n742), .d(new_n741), .O(new_n1248));
  aoi21 g0863(.a(new_n1248), .b(new_n403), .c(new_n401), .O(\grant79 ));
  nand4 g0864(.a(new_n401), .b(new_n402), .c(new_n742), .d(new_n741), .O(new_n1250));
  aoi21 g0865(.a(\req78 ), .b(new_n742), .c(\req79 ), .O(new_n1251));
  oai21 g0866(.a(new_n1250), .b(new_n1245), .c(new_n1251), .O(new_n1252));
  aoi21 g0867(.a(new_n1252), .b(new_n747), .c(new_n749), .O(\grant80 ));
  nand2 g0868(.a(new_n1252), .b(new_n747), .O(new_n1254));
  nor2  g0869(.a(\req80 ), .b(\priority81 ), .O(new_n1255));
  nand2 g0870(.a(new_n1255), .b(new_n1254), .O(new_n1256));
  aoi21 g0871(.a(new_n1256), .b(new_n748), .c(new_n750), .O(\grant81 ));
  nor2  g0872(.a(\req81 ), .b(\priority82 ), .O(new_n1258));
  nand3 g0873(.a(new_n1258), .b(new_n1255), .c(new_n1254), .O(new_n1259));
  aoi21 g0874(.a(new_n750), .b(\priority81 ), .c(\priority82 ), .O(new_n1260));
  aoi21 g0875(.a(new_n1260), .b(new_n1259), .c(new_n758), .O(\grant82 ));
  aoi21 g0876(.a(new_n1260), .b(new_n1259), .c(\req82 ), .O(new_n1262));
  inv1  g0877(.a(new_n1262), .O(new_n1263));
  aoi21 g0878(.a(new_n1263), .b(new_n756), .c(new_n399), .O(\grant83 ));
  inv1  g0879(.a(\req84 ), .O(new_n1265));
  nand4 g0880(.a(new_n1262), .b(new_n399), .c(new_n757), .d(new_n756), .O(new_n1266));
  aoi21 g0881(.a(new_n1266), .b(new_n400), .c(new_n1265), .O(\grant84 ));
  nand4 g0882(.a(new_n1265), .b(new_n399), .c(new_n757), .d(new_n756), .O(new_n1268));
  aoi21 g0883(.a(\req83 ), .b(new_n757), .c(\req84 ), .O(new_n1269));
  oai21 g0884(.a(new_n1268), .b(new_n1262), .c(new_n1269), .O(new_n1270));
  aoi21 g0885(.a(new_n1270), .b(new_n763), .c(new_n765), .O(\grant85 ));
  nand2 g0886(.a(new_n1270), .b(new_n763), .O(new_n1272));
  nor2  g0887(.a(\req85 ), .b(\priority86 ), .O(new_n1273));
  nand2 g0888(.a(new_n1273), .b(new_n1272), .O(new_n1274));
  aoi21 g0889(.a(new_n1274), .b(new_n764), .c(new_n766), .O(\grant86 ));
  nor2  g0890(.a(\req86 ), .b(\priority87 ), .O(new_n1276));
  nand3 g0891(.a(new_n1276), .b(new_n1273), .c(new_n1272), .O(new_n1277));
  aoi21 g0892(.a(new_n766), .b(\priority86 ), .c(\priority87 ), .O(new_n1278));
  aoi21 g0893(.a(new_n1278), .b(new_n1277), .c(new_n772), .O(\grant87 ));
  aoi21 g0894(.a(new_n1278), .b(new_n1277), .c(\req87 ), .O(new_n1280));
  inv1  g0895(.a(new_n1280), .O(new_n1281));
  aoi21 g0896(.a(new_n1281), .b(new_n770), .c(new_n395), .O(\grant88 ));
  nand4 g0897(.a(new_n1280), .b(new_n395), .c(new_n771), .d(new_n770), .O(new_n1283));
  aoi21 g0898(.a(new_n1283), .b(new_n396), .c(new_n394), .O(\grant89 ));
  nand4 g0899(.a(new_n394), .b(new_n395), .c(new_n771), .d(new_n770), .O(new_n1285));
  aoi21 g0900(.a(\req88 ), .b(new_n771), .c(\req89 ), .O(new_n1286));
  oai21 g0901(.a(new_n1285), .b(new_n1280), .c(new_n1286), .O(new_n1287));
  aoi21 g0902(.a(new_n1287), .b(new_n776), .c(new_n778), .O(\grant90 ));
  nand2 g0903(.a(new_n1287), .b(new_n776), .O(new_n1289));
  nor2  g0904(.a(\req90 ), .b(\priority91 ), .O(new_n1290));
  nand2 g0905(.a(new_n1290), .b(new_n1289), .O(new_n1291));
  aoi21 g0906(.a(new_n1291), .b(new_n777), .c(new_n779), .O(\grant91 ));
  inv1  g0907(.a(\req92 ), .O(new_n1293));
  nor2  g0908(.a(\req91 ), .b(\priority92 ), .O(new_n1294));
  nand3 g0909(.a(new_n1294), .b(new_n1290), .c(new_n1289), .O(new_n1295));
  aoi21 g0910(.a(new_n779), .b(\priority91 ), .c(\priority92 ), .O(new_n1296));
  aoi21 g0911(.a(new_n1296), .b(new_n1295), .c(new_n1293), .O(\grant92 ));
  nand2 g0912(.a(new_n1296), .b(new_n1295), .O(new_n1298));
  aoi21 g0913(.a(new_n1298), .b(new_n1293), .c(\priority93 ), .O(new_n1299));
  nor2  g0914(.a(new_n1299), .b(new_n392), .O(\grant93 ));
  inv1  g0915(.a(\req94 ), .O(new_n1301));
  nand3 g0916(.a(new_n1298), .b(new_n786), .c(new_n785), .O(new_n1302));
  aoi21 g0917(.a(new_n1302), .b(new_n393), .c(new_n1301), .O(\grant94 ));
  nand2 g0918(.a(new_n1302), .b(new_n393), .O(new_n1304));
  nor2  g0919(.a(\req94 ), .b(\priority95 ), .O(new_n1305));
  nand2 g0920(.a(new_n1305), .b(new_n1304), .O(new_n1306));
  aoi21 g0921(.a(new_n1306), .b(new_n791), .c(new_n793), .O(\grant95 ));
  nor2  g0922(.a(\req95 ), .b(\priority96 ), .O(new_n1308));
  nand3 g0923(.a(new_n1308), .b(new_n1305), .c(new_n1304), .O(new_n1309));
  aoi21 g0924(.a(new_n793), .b(\priority95 ), .c(\priority96 ), .O(new_n1310));
  aoi21 g0925(.a(new_n1310), .b(new_n1309), .c(new_n794), .O(\grant96 ));
  inv1  g0926(.a(\req97 ), .O(new_n1312));
  aoi21 g0927(.a(new_n1310), .b(new_n1309), .c(\req96 ), .O(new_n1313));
  inv1  g0928(.a(new_n1313), .O(new_n1314));
  aoi21 g0929(.a(new_n1314), .b(new_n391), .c(new_n1312), .O(\grant97 ));
  inv1  g0930(.a(\req98 ), .O(new_n1316));
  nand4 g0931(.a(new_n1313), .b(new_n1312), .c(new_n798), .d(new_n391), .O(new_n1317));
  aoi21 g0932(.a(new_n1312), .b(\priority97 ), .c(\priority98 ), .O(new_n1318));
  aoi21 g0933(.a(new_n1318), .b(new_n1317), .c(new_n1316), .O(\grant98 ));
  nand3 g0934(.a(new_n800), .b(new_n798), .c(new_n391), .O(new_n1320));
  aoi21 g0935(.a(\req97 ), .b(new_n798), .c(\req98 ), .O(new_n1321));
  oai21 g0936(.a(new_n1320), .b(new_n1313), .c(new_n1321), .O(new_n1322));
  aoi21 g0937(.a(new_n1322), .b(new_n799), .c(new_n390), .O(\grant99 ));
  nand2 g0938(.a(new_n1322), .b(new_n799), .O(new_n1324));
  nor2  g0939(.a(\req99 ), .b(\priority100 ), .O(new_n1325));
  nand2 g0940(.a(new_n1325), .b(new_n1324), .O(new_n1326));
  aoi21 g0941(.a(new_n1326), .b(new_n805), .c(new_n807), .O(\grant100 ));
  nand4 g0942(.a(new_n1325), .b(new_n1324), .c(new_n807), .d(new_n806), .O(new_n1328));
  aoi21 g0943(.a(new_n807), .b(\priority100 ), .c(\priority101 ), .O(new_n1329));
  aoi21 g0944(.a(new_n1329), .b(new_n1328), .c(new_n808), .O(\grant101 ));
  inv1  g0945(.a(\priority102 ), .O(new_n1331));
  inv1  g0946(.a(\req102 ), .O(new_n1332));
  nor3  g0947(.a(\req100 ), .b(\req99 ), .c(\priority100 ), .O(new_n1333));
  nand3 g0948(.a(new_n1333), .b(new_n1322), .c(new_n799), .O(new_n1334));
  aoi21 g0949(.a(\req99 ), .b(new_n805), .c(\req100 ), .O(new_n1335));
  nand2 g0950(.a(new_n1335), .b(new_n1334), .O(new_n1336));
  nand2 g0951(.a(new_n1336), .b(new_n806), .O(new_n1337));
  nor2  g0952(.a(\req101 ), .b(\priority102 ), .O(new_n1338));
  nand2 g0953(.a(new_n1338), .b(new_n1337), .O(new_n1339));
  aoi21 g0954(.a(new_n1339), .b(new_n1331), .c(new_n1332), .O(\grant102 ));
  inv1  g0955(.a(\req103 ), .O(new_n1341));
  nand3 g0956(.a(new_n1338), .b(new_n1337), .c(new_n833), .O(new_n1342));
  aoi21 g0957(.a(new_n1332), .b(\priority102 ), .c(\priority103 ), .O(new_n1343));
  aoi21 g0958(.a(new_n1343), .b(new_n1342), .c(new_n1341), .O(\grant103 ));
  inv1  g0959(.a(\req104 ), .O(new_n1345));
  aoi21 g0960(.a(new_n1343), .b(new_n1342), .c(\req103 ), .O(new_n1346));
  inv1  g0961(.a(new_n1346), .O(new_n1347));
  aoi21 g0962(.a(new_n1347), .b(new_n817), .c(new_n1345), .O(\grant104 ));
  inv1  g0963(.a(\priority105 ), .O(new_n1349));
  nand4 g0964(.a(new_n1346), .b(new_n1345), .c(new_n1349), .d(new_n817), .O(new_n1350));
  aoi21 g0965(.a(new_n1345), .b(\priority104 ), .c(\priority105 ), .O(new_n1351));
  aoi21 g0966(.a(new_n1351), .b(new_n1350), .c(new_n821), .O(\grant105 ));
  inv1  g0967(.a(\priority106 ), .O(new_n1353));
  nand4 g0968(.a(new_n821), .b(new_n1345), .c(new_n1349), .d(new_n817), .O(new_n1354));
  aoi21 g0969(.a(\req104 ), .b(new_n1349), .c(\req105 ), .O(new_n1355));
  oai21 g0970(.a(new_n1354), .b(new_n1346), .c(new_n1355), .O(new_n1356));
  aoi21 g0971(.a(new_n1356), .b(new_n1353), .c(new_n816), .O(\grant106 ));
  inv1  g0972(.a(\req107 ), .O(new_n1358));
  nand2 g0973(.a(new_n1356), .b(new_n1353), .O(new_n1359));
  nor2  g0974(.a(\req106 ), .b(\priority107 ), .O(new_n1360));
  nand2 g0975(.a(new_n1360), .b(new_n1359), .O(new_n1361));
  aoi21 g0976(.a(new_n1361), .b(new_n814), .c(new_n1358), .O(\grant107 ));
  inv1  g0977(.a(\req108 ), .O(new_n1363));
  nor2  g0978(.a(\req107 ), .b(\priority108 ), .O(new_n1364));
  nand3 g0979(.a(new_n1364), .b(new_n1360), .c(new_n1359), .O(new_n1365));
  aoi21 g0980(.a(new_n1358), .b(\priority107 ), .c(\priority108 ), .O(new_n1366));
  aoi21 g0981(.a(new_n1366), .b(new_n1365), .c(new_n1363), .O(\grant108 ));
  inv1  g0982(.a(\req109 ), .O(new_n1368));
  inv1  g0983(.a(new_n828), .O(new_n1369));
  nand2 g0984(.a(new_n1329), .b(new_n1328), .O(new_n1370));
  nand2 g0985(.a(new_n1370), .b(new_n808), .O(new_n1371));
  nor4  g0986(.a(new_n831), .b(\req102 ), .c(\priority103 ), .d(\priority102 ), .O(new_n1372));
  oai21 g0987(.a(new_n1332), .b(\priority103 ), .c(new_n832), .O(new_n1373));
  aoi21 g0988(.a(new_n1372), .b(new_n1371), .c(new_n1373), .O(new_n1374));
  nor2  g0989(.a(new_n1374), .b(new_n1369), .O(new_n1375));
  nor2  g0990(.a(new_n1375), .b(new_n1368), .O(\grant109 ));
  nor2  g0991(.a(\req109 ), .b(\priority110 ), .O(new_n1377));
  oai21 g0992(.a(new_n1374), .b(new_n1369), .c(new_n1377), .O(new_n1378));
  aoi21 g0993(.a(new_n1378), .b(new_n841), .c(new_n843), .O(\grant110 ));
  nand4 g0994(.a(new_n840), .b(new_n843), .c(new_n842), .d(new_n841), .O(new_n1380));
  aoi21 g0995(.a(new_n843), .b(\priority110 ), .c(\priority111 ), .O(new_n1381));
  aoi21 g0996(.a(new_n1381), .b(new_n1380), .c(new_n844), .O(\grant111 ));
  nand2 g0997(.a(new_n847), .b(new_n389), .O(new_n1383));
  inv1  g0998(.a(new_n1383), .O(new_n1384));
  nor2  g0999(.a(new_n1384), .b(new_n450), .O(\grant112 ));
  nor3  g1000(.a(new_n1384), .b(\req112 ), .c(\priority113 ), .O(new_n1386));
  inv1  g1001(.a(new_n1386), .O(new_n1387));
  aoi21 g1002(.a(new_n1387), .b(new_n449), .c(new_n447), .O(\grant113 ));
  inv1  g1003(.a(\req114 ), .O(new_n1389));
  nand2 g1004(.a(new_n1386), .b(new_n451), .O(new_n1390));
  aoi21 g1005(.a(new_n1390), .b(new_n448), .c(new_n1389), .O(\grant114 ));
  aoi21 g1006(.a(new_n852), .b(new_n1389), .c(\priority115 ), .O(new_n1392));
  nor2  g1007(.a(new_n1392), .b(new_n856), .O(\grant115 ));
  aoi21 g1008(.a(new_n857), .b(new_n855), .c(new_n437), .O(\grant116 ));
  aoi21 g1009(.a(new_n858), .b(new_n437), .c(\priority117 ), .O(new_n1395));
  nor2  g1010(.a(new_n1395), .b(new_n435), .O(\grant117 ));
  aoi21 g1011(.a(new_n862), .b(new_n861), .c(new_n457), .O(\grant118 ));
  inv1  g1012(.a(\req119 ), .O(new_n1398));
  inv1  g1013(.a(new_n863), .O(new_n1399));
  aoi21 g1014(.a(new_n1399), .b(new_n456), .c(new_n1398), .O(\grant119 ));
  inv1  g1015(.a(\req120 ), .O(new_n1401));
  nand4 g1016(.a(new_n863), .b(new_n1398), .c(new_n864), .d(new_n456), .O(new_n1402));
  aoi21 g1017(.a(new_n1398), .b(\priority119 ), .c(\priority120 ), .O(new_n1403));
  aoi21 g1018(.a(new_n1403), .b(new_n1402), .c(new_n1401), .O(\grant120 ));
  inv1  g1019(.a(new_n868), .O(new_n1405));
  nor2  g1020(.a(new_n1405), .b(new_n429), .O(\grant121 ));
  nor3  g1021(.a(new_n1405), .b(\req121 ), .c(\priority122 ), .O(new_n1407));
  inv1  g1022(.a(new_n1407), .O(new_n1408));
  aoi21 g1023(.a(new_n1408), .b(new_n869), .c(new_n430), .O(\grant122 ));
  nand3 g1024(.a(new_n1407), .b(new_n430), .c(new_n468), .O(new_n1410));
  aoi21 g1025(.a(new_n430), .b(\priority122 ), .c(\priority123 ), .O(new_n1411));
  aoi21 g1026(.a(new_n1411), .b(new_n1410), .c(new_n870), .O(\grant123 ));
  aoi21 g1027(.a(new_n878), .b(new_n469), .c(new_n879), .O(\grant124 ));
  inv1  g1028(.a(new_n878), .O(new_n1414));
  nand4 g1029(.a(new_n1414), .b(new_n879), .c(new_n473), .d(new_n469), .O(new_n1415));
  aoi21 g1030(.a(new_n879), .b(\priority124 ), .c(\priority125 ), .O(new_n1416));
  aoi21 g1031(.a(new_n1416), .b(new_n1415), .c(new_n475), .O(\grant125 ));
  nor2  g1032(.a(new_n883), .b(\priority126 ), .O(new_n1418));
  nor2  g1033(.a(new_n1418), .b(new_n476), .O(\grant126 ));
  inv1  g1034(.a(\priority127 ), .O(new_n1420));
  aoi21 g1035(.a(new_n885), .b(new_n1420), .c(new_n888), .O(\grant127 ));
  nand3 g1036(.a(new_n844), .b(new_n843), .c(new_n1368), .O(new_n1422));
  nand4 g1037(.a(new_n1332), .b(new_n1316), .c(new_n1312), .d(new_n794), .O(new_n1423));
  nand4 g1038(.a(new_n793), .b(new_n1301), .c(new_n392), .d(new_n1293), .O(new_n1424));
  nor3  g1039(.a(new_n1424), .b(new_n1423), .c(new_n1422), .O(new_n1425));
  nand3 g1040(.a(new_n1425), .b(new_n589), .c(new_n416), .O(new_n1426));
  nand4 g1041(.a(new_n512), .b(new_n505), .c(new_n497), .d(new_n489), .O(new_n1427));
  inv1  g1042(.a(new_n1427), .O(new_n1428));
  nand4 g1043(.a(new_n1428), .b(new_n832), .c(new_n434), .d(new_n446), .O(new_n1429));
  nand4 g1044(.a(new_n750), .b(new_n749), .c(new_n402), .d(new_n737), .O(new_n1430));
  nand4 g1045(.a(new_n689), .b(new_n688), .c(new_n680), .d(new_n679), .O(new_n1431));
  nor2  g1046(.a(new_n1431), .b(new_n1430), .O(new_n1432));
  nand4 g1047(.a(new_n779), .b(new_n394), .c(new_n395), .d(new_n772), .O(new_n1433));
  nand4 g1048(.a(new_n765), .b(new_n1265), .c(new_n399), .d(new_n758), .O(new_n1434));
  nor2  g1049(.a(new_n1434), .b(new_n1433), .O(new_n1435));
  nand2 g1050(.a(new_n1435), .b(new_n1432), .O(new_n1436));
  nand4 g1051(.a(new_n630), .b(new_n629), .c(new_n621), .d(new_n620), .O(new_n1437));
  nand4 g1052(.a(new_n1071), .b(new_n603), .c(new_n594), .d(new_n426), .O(new_n1438));
  nor2  g1053(.a(new_n1438), .b(new_n1437), .O(new_n1439));
  nand3 g1054(.a(new_n1147), .b(new_n664), .c(new_n663), .O(new_n1440));
  nand4 g1055(.a(new_n655), .b(new_n1122), .c(new_n645), .d(new_n637), .O(new_n1441));
  nor2  g1056(.a(new_n1441), .b(new_n1440), .O(new_n1442));
  nand2 g1057(.a(new_n1442), .b(new_n1439), .O(new_n1443));
  nor4  g1058(.a(new_n1443), .b(new_n1436), .c(new_n1429), .d(new_n1426), .O(new_n1444));
  nor2  g1059(.a(\req3 ), .b(\req1 ), .O(new_n1445));
  nor2  g1060(.a(\req79 ), .b(\req77 ), .O(new_n1446));
  nand4 g1061(.a(new_n1446), .b(new_n1445), .c(new_n736), .d(new_n421), .O(new_n1447));
  inv1  g1062(.a(new_n1447), .O(new_n1448));
  nor2  g1063(.a(\req36 ), .b(\req34 ), .O(new_n1449));
  nand4 g1064(.a(new_n1449), .b(new_n483), .c(new_n595), .d(new_n914), .O(new_n1450));
  nand4 g1065(.a(new_n778), .b(new_n766), .c(new_n1228), .d(new_n1160), .O(new_n1451));
  nand4 g1066(.a(new_n671), .b(new_n654), .c(new_n646), .d(new_n612), .O(new_n1452));
  nor3  g1067(.a(\req125 ), .b(\req113 ), .c(\req5 ), .O(new_n1453));
  nor2  g1068(.a(\req112 ), .b(\req101 ), .O(new_n1454));
  nand4 g1069(.a(new_n1454), .b(new_n1453), .c(new_n807), .d(new_n390), .O(new_n1455));
  nor4  g1070(.a(new_n1455), .b(new_n1452), .c(new_n1451), .d(new_n1450), .O(new_n1456));
  inv1  g1071(.a(new_n1444), .O(new_n1457));
  nor2  g1072(.a(new_n1447), .b(new_n1457), .O(new_n1458));
  nand2 g1073(.a(new_n1456), .b(new_n521), .O(new_n1459));
  inv1  g1074(.a(new_n1459), .O(new_n1460));
  inv1  g1075(.a(new_n521), .O(new_n1461));
  nand3 g1076(.a(new_n1456), .b(new_n1461), .c(\req44 ), .O(new_n1462));
  inv1  g1077(.a(new_n1462), .O(new_n1463));
  oai21 g1078(.a(new_n1463), .b(new_n1460), .c(new_n1458), .O(new_n1464));
  nand4 g1079(.a(new_n1464), .b(new_n1456), .c(new_n1448), .d(new_n1444), .O(anyGrant));
endmodule


